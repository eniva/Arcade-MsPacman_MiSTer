library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"3E",X"3F",X"ED",X"47",X"C3",X"0B",X"23",X"77",X"23",X"10",X"FC",X"C9",X"C3",X"0E",X"07",
		X"85",X"6F",X"3E",X"00",X"8C",X"67",X"7E",X"C9",X"78",X"87",X"D7",X"5F",X"23",X"56",X"EB",X"C9",
		X"E1",X"87",X"D7",X"5F",X"23",X"56",X"EB",X"E9",X"E1",X"46",X"23",X"4E",X"23",X"E5",X"18",X"12",
		X"11",X"90",X"4C",X"06",X"10",X"C3",X"51",X"00",X"AF",X"32",X"00",X"50",X"32",X"07",X"50",X"C3",
		X"38",X"00",X"2A",X"80",X"4C",X"70",X"2C",X"71",X"2C",X"20",X"02",X"2E",X"C0",X"22",X"80",X"4C",
		X"C9",X"1A",X"A7",X"28",X"06",X"1C",X"1C",X"1C",X"10",X"F7",X"C9",X"E1",X"06",X"03",X"7E",X"12",
		X"23",X"1C",X"10",X"FA",X"E9",X"C3",X"2D",X"20",X"00",X"01",X"02",X"03",X"04",X"05",X"06",X"07",
		X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"12",X"13",X"14",X"01",X"03",X"04",
		X"06",X"07",X"08",X"09",X"0A",X"0B",X"0C",X"0D",X"0E",X"0F",X"10",X"11",X"14",X"F5",X"32",X"C0",
		X"50",X"AF",X"32",X"00",X"50",X"F3",X"C5",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"21",X"8C",X"4E",
		X"11",X"50",X"50",X"01",X"10",X"00",X"ED",X"B0",X"3A",X"CC",X"4E",X"A7",X"3A",X"CF",X"4E",X"20",
		X"03",X"3A",X"9F",X"4E",X"32",X"45",X"50",X"3A",X"DC",X"4E",X"A7",X"3A",X"DF",X"4E",X"20",X"03",
		X"3A",X"AF",X"4E",X"32",X"4A",X"50",X"3A",X"EC",X"4E",X"A7",X"3A",X"EF",X"4E",X"20",X"03",X"3A",
		X"BF",X"4E",X"32",X"4F",X"50",X"21",X"02",X"4C",X"11",X"22",X"4C",X"01",X"1C",X"00",X"ED",X"B0",
		X"DD",X"21",X"20",X"4C",X"DD",X"7E",X"02",X"07",X"07",X"DD",X"77",X"02",X"DD",X"7E",X"04",X"07",
		X"07",X"DD",X"77",X"04",X"DD",X"7E",X"06",X"07",X"07",X"DD",X"77",X"06",X"DD",X"7E",X"08",X"07",
		X"07",X"DD",X"77",X"08",X"DD",X"7E",X"0A",X"07",X"07",X"DD",X"77",X"0A",X"DD",X"7E",X"0C",X"07",
		X"07",X"DD",X"77",X"0C",X"3A",X"D1",X"4D",X"FE",X"01",X"20",X"38",X"DD",X"21",X"20",X"4C",X"3A",
		X"A4",X"4D",X"87",X"5F",X"16",X"00",X"DD",X"19",X"2A",X"24",X"4C",X"ED",X"5B",X"34",X"4C",X"DD",
		X"7E",X"00",X"32",X"24",X"4C",X"DD",X"7E",X"01",X"32",X"25",X"4C",X"DD",X"7E",X"10",X"32",X"34",
		X"4C",X"DD",X"7E",X"11",X"32",X"35",X"4C",X"DD",X"75",X"00",X"DD",X"74",X"01",X"DD",X"73",X"10",
		X"DD",X"72",X"11",X"3A",X"A6",X"4D",X"A7",X"CA",X"76",X"01",X"ED",X"4B",X"22",X"4C",X"ED",X"5B",
		X"32",X"4C",X"2A",X"2A",X"4C",X"22",X"22",X"4C",X"2A",X"3A",X"4C",X"22",X"32",X"4C",X"ED",X"43",
		X"2A",X"4C",X"ED",X"53",X"3A",X"4C",X"21",X"22",X"4C",X"11",X"F2",X"4F",X"01",X"0C",X"00",X"ED",
		X"B0",X"21",X"32",X"4C",X"11",X"62",X"50",X"01",X"0C",X"00",X"ED",X"B0",X"CD",X"DC",X"01",X"CD",
		X"21",X"02",X"CD",X"C8",X"03",X"3A",X"00",X"4E",X"A7",X"28",X"12",X"CD",X"9D",X"03",X"CD",X"90",
		X"14",X"CD",X"1F",X"14",X"CD",X"67",X"02",X"CD",X"AD",X"02",X"CD",X"FD",X"02",X"3A",X"00",X"4E",
		X"3D",X"20",X"06",X"32",X"AC",X"4E",X"32",X"BC",X"4E",X"CD",X"0C",X"2D",X"CD",X"C1",X"2C",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"D1",X"C1",X"3A",X"00",X"4E",X"A7",X"28",X"08",X"3A",X"40",X"50",X"E6",
		X"10",X"CA",X"00",X"00",X"3E",X"01",X"32",X"00",X"50",X"FB",X"F1",X"C9",X"21",X"84",X"4C",X"34",
		X"23",X"35",X"23",X"11",X"19",X"02",X"01",X"01",X"04",X"34",X"7E",X"E6",X"0F",X"EB",X"BE",X"20",
		X"13",X"0C",X"1A",X"C6",X"10",X"E6",X"F0",X"12",X"23",X"BE",X"20",X"08",X"0C",X"EB",X"36",X"00",
		X"23",X"13",X"10",X"E5",X"21",X"8A",X"4C",X"71",X"2C",X"7E",X"87",X"87",X"86",X"3C",X"77",X"2C",
		X"7E",X"87",X"86",X"87",X"87",X"86",X"3C",X"77",X"C9",X"06",X"A0",X"0A",X"60",X"0A",X"60",X"0A",
		X"A0",X"21",X"90",X"4C",X"3A",X"8A",X"4C",X"4F",X"06",X"10",X"7E",X"A7",X"28",X"2F",X"E6",X"C0",
		X"07",X"07",X"B9",X"30",X"28",X"35",X"7E",X"E6",X"3F",X"20",X"22",X"77",X"C5",X"E5",X"2C",X"7E",
		X"2C",X"46",X"21",X"5B",X"02",X"E5",X"E7",X"94",X"08",X"A3",X"06",X"8E",X"05",X"72",X"12",X"00",
		X"10",X"0B",X"10",X"63",X"02",X"2B",X"21",X"F0",X"21",X"B9",X"22",X"E1",X"C1",X"2C",X"2C",X"2C",
		X"10",X"C8",X"C9",X"EF",X"1C",X"86",X"C9",X"3A",X"6E",X"4E",X"FE",X"99",X"17",X"32",X"06",X"50",
		X"1F",X"D0",X"3A",X"00",X"50",X"47",X"CB",X"00",X"3A",X"66",X"4E",X"17",X"E6",X"0F",X"32",X"66",
		X"4E",X"D6",X"0C",X"CC",X"DF",X"02",X"CB",X"00",X"3A",X"67",X"4E",X"17",X"E6",X"0F",X"32",X"67",
		X"4E",X"D6",X"0C",X"C2",X"9A",X"02",X"21",X"69",X"4E",X"34",X"CB",X"00",X"3A",X"68",X"4E",X"17",
		X"E6",X"0F",X"32",X"68",X"4E",X"D6",X"0C",X"C0",X"21",X"69",X"4E",X"34",X"C9",X"3A",X"69",X"4E",
		X"A7",X"C8",X"47",X"3A",X"6A",X"4E",X"5F",X"FE",X"00",X"C2",X"C4",X"02",X"3E",X"01",X"32",X"07",
		X"50",X"CD",X"DF",X"02",X"7B",X"FE",X"08",X"C2",X"CE",X"02",X"AF",X"32",X"07",X"50",X"1C",X"7B",
		X"32",X"6A",X"4E",X"D6",X"10",X"C0",X"32",X"6A",X"4E",X"05",X"78",X"32",X"69",X"4E",X"C9",X"3A",
		X"6B",X"4E",X"21",X"6C",X"4E",X"34",X"96",X"C0",X"77",X"3A",X"6D",X"4E",X"21",X"6E",X"4E",X"86",
		X"27",X"D2",X"F6",X"02",X"3E",X"99",X"77",X"21",X"9C",X"4E",X"CB",X"CE",X"C9",X"21",X"CE",X"4D",
		X"34",X"7E",X"E6",X"0F",X"20",X"1F",X"7E",X"0F",X"0F",X"0F",X"0F",X"47",X"3A",X"D6",X"4D",X"2F",
		X"B0",X"4F",X"3A",X"6E",X"4E",X"D6",X"01",X"30",X"02",X"AF",X"4F",X"28",X"01",X"79",X"32",X"05",
		X"50",X"79",X"32",X"04",X"50",X"DD",X"21",X"D8",X"43",X"FD",X"21",X"C5",X"43",X"3A",X"00",X"4E",
		X"FE",X"03",X"CA",X"44",X"03",X"3A",X"03",X"4E",X"FE",X"02",X"D2",X"44",X"03",X"CD",X"69",X"03",
		X"CD",X"76",X"03",X"C9",X"3A",X"09",X"4E",X"A7",X"3A",X"CE",X"4D",X"C2",X"59",X"03",X"CB",X"67",
		X"CC",X"69",X"03",X"C4",X"83",X"03",X"C3",X"61",X"03",X"CB",X"67",X"CC",X"76",X"03",X"C4",X"90",
		X"03",X"3A",X"70",X"4E",X"A7",X"CC",X"90",X"03",X"C9",X"DD",X"36",X"00",X"50",X"DD",X"36",X"01",
		X"55",X"DD",X"36",X"02",X"31",X"C9",X"FD",X"36",X"00",X"50",X"FD",X"36",X"01",X"55",X"FD",X"36",
		X"02",X"32",X"C9",X"DD",X"36",X"00",X"40",X"DD",X"36",X"01",X"40",X"DD",X"36",X"02",X"40",X"C9",
		X"FD",X"36",X"00",X"40",X"FD",X"36",X"01",X"40",X"FD",X"36",X"02",X"40",X"C9",X"3A",X"06",X"4E",
		X"D6",X"05",X"D8",X"2A",X"08",X"4D",X"06",X"08",X"0E",X"10",X"7D",X"32",X"06",X"4D",X"32",X"D2",
		X"4D",X"91",X"32",X"02",X"4D",X"32",X"04",X"4D",X"7C",X"80",X"32",X"03",X"4D",X"32",X"07",X"4D",
		X"91",X"32",X"05",X"4D",X"32",X"D3",X"4D",X"C9",X"3A",X"00",X"4E",X"E7",X"D4",X"03",X"FE",X"03",
		X"E5",X"05",X"BE",X"06",X"3A",X"01",X"4E",X"E7",X"DC",X"03",X"0C",X"00",X"EF",X"00",X"00",X"EF",
		X"06",X"00",X"EF",X"01",X"00",X"EF",X"14",X"00",X"EF",X"18",X"00",X"EF",X"04",X"00",X"EF",X"1E",
		X"00",X"EF",X"07",X"00",X"21",X"01",X"4E",X"34",X"21",X"01",X"50",X"36",X"01",X"C9",X"CD",X"A1",
		X"2B",X"3A",X"6E",X"4E",X"A7",X"28",X"0C",X"AF",X"32",X"04",X"4E",X"32",X"02",X"4E",X"21",X"00",
		X"4E",X"34",X"C9",X"3A",X"02",X"4E",X"E7",X"5F",X"04",X"0C",X"00",X"71",X"04",X"0C",X"00",X"7F",
		X"04",X"0C",X"00",X"85",X"04",X"0C",X"00",X"8B",X"04",X"0C",X"00",X"99",X"04",X"0C",X"00",X"9F",
		X"04",X"0C",X"00",X"A5",X"04",X"0C",X"00",X"B3",X"04",X"0C",X"00",X"B9",X"04",X"0C",X"00",X"BF",
		X"04",X"0C",X"00",X"CD",X"04",X"0C",X"00",X"D3",X"04",X"0C",X"00",X"D8",X"04",X"0C",X"00",X"E0",
		X"04",X"0C",X"00",X"1C",X"05",X"4B",X"05",X"56",X"05",X"61",X"05",X"6C",X"05",X"7C",X"05",X"EF",
		X"00",X"01",X"EF",X"01",X"00",X"EF",X"04",X"00",X"EF",X"1E",X"00",X"0E",X"0C",X"CD",X"85",X"05",
		X"C9",X"21",X"04",X"43",X"3E",X"01",X"CD",X"BF",X"05",X"0E",X"0C",X"CD",X"85",X"05",X"C9",X"0E",
		X"14",X"CD",X"93",X"05",X"C9",X"0E",X"0D",X"CD",X"93",X"05",X"C9",X"21",X"07",X"43",X"3E",X"03",
		X"CD",X"BF",X"05",X"0E",X"0C",X"CD",X"85",X"05",X"C9",X"0E",X"16",X"CD",X"93",X"05",X"C9",X"0E",
		X"0F",X"CD",X"93",X"05",X"C9",X"21",X"0A",X"43",X"3E",X"05",X"CD",X"BF",X"05",X"0E",X"0C",X"CD",
		X"85",X"05",X"C9",X"0E",X"33",X"CD",X"93",X"05",X"C9",X"0E",X"2F",X"CD",X"93",X"05",X"C9",X"21",
		X"0D",X"43",X"3E",X"07",X"CD",X"BF",X"05",X"0E",X"0C",X"CD",X"85",X"05",X"C9",X"0E",X"35",X"CD",
		X"93",X"05",X"C9",X"0E",X"31",X"C3",X"80",X"05",X"EF",X"1C",X"11",X"0E",X"12",X"C3",X"85",X"05",
		X"0E",X"13",X"CD",X"85",X"05",X"CD",X"79",X"08",X"35",X"EF",X"11",X"00",X"EF",X"05",X"01",X"EF",
		X"10",X"14",X"EF",X"04",X"01",X"3E",X"01",X"32",X"14",X"4E",X"AF",X"32",X"70",X"4E",X"32",X"15",
		X"4E",X"21",X"32",X"43",X"36",X"14",X"3E",X"FC",X"11",X"20",X"00",X"06",X"1C",X"DD",X"21",X"40",
		X"40",X"DD",X"77",X"11",X"DD",X"77",X"13",X"DD",X"19",X"10",X"F6",X"C9",X"21",X"A0",X"4D",X"06",
		X"21",X"3A",X"3A",X"4D",X"90",X"20",X"05",X"36",X"01",X"C3",X"8E",X"05",X"CD",X"17",X"10",X"CD",
		X"17",X"10",X"CD",X"23",X"0E",X"CD",X"0D",X"0C",X"CD",X"D6",X"0B",X"CD",X"A5",X"05",X"CD",X"FE",
		X"1E",X"CD",X"25",X"1F",X"CD",X"4C",X"1F",X"CD",X"73",X"1F",X"C9",X"21",X"A1",X"4D",X"06",X"20",
		X"3A",X"32",X"4D",X"C3",X"24",X"05",X"21",X"A2",X"4D",X"06",X"22",X"3A",X"32",X"4D",X"C3",X"24",
		X"05",X"21",X"A3",X"4D",X"06",X"24",X"3A",X"32",X"4D",X"C3",X"24",X"05",X"3A",X"D0",X"4D",X"47",
		X"3A",X"D1",X"4D",X"80",X"FE",X"06",X"CA",X"8E",X"05",X"C3",X"2C",X"05",X"CD",X"BE",X"06",X"C9",
		X"3A",X"75",X"4E",X"81",X"4F",X"06",X"1C",X"CD",X"42",X"00",X"F7",X"4A",X"02",X"00",X"21",X"02",
		X"4E",X"34",X"C9",X"3A",X"75",X"4E",X"81",X"4F",X"06",X"1C",X"CD",X"42",X"00",X"F7",X"45",X"02",
		X"00",X"CD",X"8E",X"05",X"C9",X"3A",X"B5",X"4D",X"A7",X"C8",X"AF",X"32",X"B5",X"4D",X"3A",X"30",
		X"4D",X"EE",X"02",X"32",X"3C",X"4D",X"47",X"21",X"FF",X"32",X"DF",X"22",X"26",X"4D",X"C9",X"36",
		X"B1",X"2C",X"36",X"B3",X"2C",X"36",X"B5",X"01",X"1E",X"00",X"09",X"36",X"B0",X"2C",X"36",X"B2",
		X"2C",X"36",X"B4",X"11",X"00",X"04",X"19",X"77",X"2D",X"77",X"2D",X"77",X"A7",X"ED",X"42",X"77",
		X"2D",X"77",X"2D",X"77",X"C9",X"3A",X"03",X"4E",X"E7",X"F3",X"05",X"1B",X"06",X"74",X"06",X"0C",
		X"00",X"A8",X"06",X"CD",X"A1",X"2B",X"EF",X"00",X"01",X"EF",X"01",X"00",X"EF",X"1C",X"07",X"EF",
		X"1C",X"0B",X"EF",X"1E",X"00",X"21",X"03",X"4E",X"34",X"3E",X"01",X"32",X"D6",X"4D",X"3A",X"71",
		X"4E",X"FE",X"FF",X"C8",X"EF",X"1C",X"0A",X"EF",X"1F",X"00",X"C9",X"CD",X"A1",X"2B",X"3A",X"6E",
		X"4E",X"FE",X"01",X"06",X"09",X"20",X"02",X"06",X"08",X"CD",X"5E",X"2C",X"3A",X"6E",X"4E",X"FE",
		X"01",X"3A",X"40",X"50",X"28",X"0C",X"CB",X"77",X"20",X"08",X"3E",X"01",X"32",X"70",X"4E",X"C3",
		X"49",X"06",X"CB",X"6F",X"C0",X"AF",X"32",X"70",X"4E",X"3A",X"6B",X"4E",X"A7",X"28",X"15",X"3A",
		X"70",X"4E",X"A7",X"3A",X"6E",X"4E",X"28",X"03",X"C6",X"99",X"27",X"C6",X"99",X"27",X"32",X"6E",
		X"4E",X"CD",X"A1",X"2B",X"21",X"03",X"4E",X"34",X"AF",X"32",X"D6",X"4D",X"3C",X"32",X"CC",X"4E",
		X"32",X"DC",X"4E",X"C9",X"EF",X"00",X"01",X"EF",X"01",X"01",X"EF",X"02",X"00",X"EF",X"12",X"00",
		X"EF",X"03",X"00",X"EF",X"1C",X"03",X"EF",X"1C",X"06",X"EF",X"18",X"00",X"EF",X"1B",X"00",X"AF",
		X"32",X"13",X"4E",X"3A",X"6F",X"4E",X"32",X"14",X"4E",X"32",X"15",X"4E",X"EF",X"1A",X"00",X"F7",
		X"57",X"01",X"00",X"21",X"03",X"4E",X"34",X"C9",X"21",X"15",X"4E",X"35",X"CD",X"6A",X"2B",X"AF",
		X"32",X"03",X"4E",X"32",X"02",X"4E",X"32",X"04",X"4E",X"21",X"00",X"4E",X"34",X"C9",X"3A",X"04",
		X"4E",X"E7",X"79",X"08",X"99",X"08",X"0C",X"00",X"CD",X"08",X"0D",X"09",X"0C",X"00",X"40",X"09",
		X"0C",X"00",X"72",X"09",X"88",X"09",X"0C",X"00",X"D2",X"09",X"D8",X"09",X"0C",X"00",X"E8",X"09",
		X"0C",X"00",X"FE",X"09",X"0C",X"00",X"02",X"0A",X"0C",X"00",X"04",X"0A",X"0C",X"00",X"06",X"0A",
		X"0C",X"00",X"08",X"0A",X"0C",X"00",X"0A",X"0A",X"0C",X"00",X"0C",X"0A",X"0C",X"00",X"0E",X"0A",
		X"0C",X"00",X"2C",X"0A",X"0C",X"00",X"7C",X"0A",X"A0",X"0A",X"0C",X"00",X"A3",X"0A",X"78",X"A7",
		X"20",X"04",X"2A",X"0A",X"4E",X"7E",X"DD",X"21",X"96",X"07",X"47",X"87",X"87",X"80",X"80",X"5F",
		X"16",X"00",X"DD",X"19",X"DD",X"7E",X"00",X"87",X"47",X"87",X"87",X"4F",X"87",X"87",X"81",X"80",
		X"5F",X"16",X"00",X"21",X"0F",X"33",X"19",X"CD",X"14",X"08",X"DD",X"7E",X"01",X"32",X"B0",X"4D",
		X"DD",X"7E",X"02",X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"43",X"08",X"19",X"CD",X"3A",X"08",
		X"DD",X"7E",X"03",X"87",X"5F",X"16",X"00",X"FD",X"21",X"4F",X"08",X"FD",X"19",X"FD",X"6E",X"00",
		X"FD",X"66",X"01",X"22",X"BB",X"4D",X"DD",X"7E",X"04",X"87",X"5F",X"16",X"00",X"FD",X"21",X"61",
		X"08",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"BD",X"4D",X"DD",X"7E",X"05",X"87",
		X"5F",X"16",X"00",X"FD",X"21",X"73",X"08",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",
		X"95",X"4D",X"CD",X"EA",X"2B",X"C9",X"03",X"01",X"01",X"00",X"02",X"00",X"04",X"01",X"02",X"01",
		X"03",X"00",X"04",X"01",X"03",X"02",X"04",X"01",X"04",X"02",X"03",X"02",X"05",X"01",X"05",X"00",
		X"03",X"02",X"06",X"02",X"05",X"01",X"03",X"03",X"03",X"02",X"05",X"02",X"03",X"03",X"06",X"02",
		X"05",X"02",X"03",X"03",X"06",X"02",X"05",X"00",X"03",X"04",X"07",X"02",X"05",X"01",X"03",X"04",
		X"03",X"02",X"05",X"02",X"03",X"04",X"06",X"02",X"05",X"02",X"03",X"05",X"07",X"02",X"05",X"00",
		X"03",X"05",X"07",X"02",X"05",X"02",X"03",X"05",X"05",X"02",X"05",X"01",X"03",X"06",X"07",X"02",
		X"05",X"02",X"03",X"06",X"07",X"02",X"05",X"02",X"03",X"06",X"08",X"02",X"05",X"02",X"03",X"06",
		X"07",X"02",X"05",X"02",X"03",X"07",X"08",X"02",X"05",X"02",X"03",X"07",X"08",X"02",X"06",X"02",
		X"03",X"07",X"08",X"02",X"11",X"46",X"4D",X"01",X"1C",X"00",X"ED",X"B0",X"01",X"0C",X"00",X"A7",
		X"ED",X"42",X"ED",X"B0",X"01",X"0C",X"00",X"A7",X"ED",X"42",X"ED",X"B0",X"01",X"0C",X"00",X"A7",
		X"ED",X"42",X"ED",X"B0",X"01",X"0E",X"00",X"ED",X"B0",X"C9",X"11",X"B8",X"4D",X"01",X"03",X"00",
		X"ED",X"B0",X"C9",X"14",X"1E",X"46",X"00",X"1E",X"3C",X"00",X"00",X"32",X"00",X"00",X"00",X"14",
		X"0A",X"1E",X"0F",X"28",X"14",X"32",X"19",X"3C",X"1E",X"50",X"28",X"64",X"32",X"78",X"3C",X"8C",
		X"46",X"C0",X"03",X"48",X"03",X"D0",X"02",X"58",X"02",X"E0",X"01",X"68",X"01",X"F0",X"00",X"78",
		X"00",X"01",X"00",X"F0",X"00",X"F0",X"00",X"B4",X"00",X"21",X"09",X"4E",X"AF",X"06",X"0B",X"CF",
		X"CD",X"C9",X"24",X"2A",X"73",X"4E",X"22",X"0A",X"4E",X"21",X"0A",X"4E",X"11",X"38",X"4E",X"01",
		X"2E",X"00",X"ED",X"B0",X"21",X"04",X"4E",X"34",X"C9",X"3A",X"00",X"4E",X"3D",X"20",X"06",X"3E",
		X"09",X"32",X"04",X"4E",X"C9",X"EF",X"11",X"00",X"EF",X"1C",X"83",X"EF",X"04",X"00",X"EF",X"05",
		X"00",X"EF",X"10",X"00",X"EF",X"1A",X"00",X"F7",X"54",X"00",X"00",X"F7",X"54",X"06",X"00",X"3A",
		X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"32",X"03",X"50",X"C3",X"94",X"08",X"3A",X"00",X"50",
		X"CB",X"67",X"C2",X"DE",X"08",X"21",X"04",X"4E",X"36",X"0E",X"EF",X"13",X"00",X"C9",X"3A",X"0E",
		X"4E",X"FE",X"F4",X"20",X"06",X"21",X"04",X"4E",X"36",X"0C",X"C9",X"CD",X"17",X"10",X"CD",X"17",
		X"10",X"CD",X"DD",X"13",X"CD",X"42",X"0C",X"CD",X"23",X"0E",X"CD",X"36",X"0E",X"CD",X"C3",X"0A",
		X"CD",X"D6",X"0B",X"CD",X"0D",X"0C",X"CD",X"6C",X"0E",X"CD",X"AD",X"0E",X"C9",X"3E",X"01",X"32",
		X"12",X"4E",X"CD",X"87",X"24",X"21",X"04",X"4E",X"34",X"3A",X"14",X"4E",X"A7",X"20",X"1F",X"3A",
		X"70",X"4E",X"A7",X"28",X"19",X"3A",X"42",X"4E",X"A7",X"28",X"13",X"3A",X"09",X"4E",X"C6",X"03",
		X"4F",X"06",X"1C",X"CD",X"42",X"00",X"EF",X"1C",X"05",X"F7",X"54",X"00",X"00",X"C9",X"34",X"C9",
		X"3A",X"70",X"4E",X"A7",X"28",X"06",X"3A",X"42",X"4E",X"A7",X"20",X"15",X"3A",X"14",X"4E",X"A7",
		X"20",X"1A",X"CD",X"A1",X"2B",X"EF",X"1C",X"05",X"F7",X"54",X"00",X"00",X"21",X"04",X"4E",X"34",
		X"C9",X"CD",X"A6",X"0A",X"3A",X"09",X"4E",X"EE",X"01",X"32",X"09",X"4E",X"3E",X"09",X"32",X"04",
		X"4E",X"C9",X"AF",X"32",X"02",X"4E",X"32",X"04",X"4E",X"32",X"70",X"4E",X"32",X"09",X"4E",X"32",
		X"03",X"50",X"3E",X"01",X"32",X"00",X"4E",X"C9",X"EF",X"00",X"01",X"EF",X"01",X"01",X"EF",X"02",
		X"00",X"EF",X"11",X"00",X"EF",X"13",X"00",X"EF",X"03",X"00",X"EF",X"04",X"00",X"EF",X"05",X"00",
		X"EF",X"10",X"00",X"EF",X"1A",X"00",X"EF",X"1C",X"06",X"3A",X"00",X"4E",X"FE",X"03",X"28",X"06",
		X"EF",X"1C",X"05",X"EF",X"1D",X"00",X"F7",X"54",X"00",X"00",X"3A",X"00",X"4E",X"3D",X"28",X"04",
		X"F7",X"54",X"06",X"00",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"32",X"03",X"50",X"C3",
		X"94",X"08",X"3E",X"03",X"32",X"04",X"4E",X"C9",X"F7",X"54",X"00",X"00",X"21",X"04",X"4E",X"34",
		X"AF",X"32",X"AC",X"4E",X"32",X"BC",X"4E",X"C9",X"0E",X"02",X"06",X"01",X"CD",X"42",X"00",X"F7",
		X"42",X"00",X"00",X"21",X"00",X"00",X"CD",X"7E",X"26",X"21",X"04",X"4E",X"34",X"C9",X"0E",X"00",
		X"18",X"E8",X"18",X"E4",X"18",X"F8",X"18",X"E0",X"18",X"F4",X"18",X"DC",X"18",X"F0",X"EF",X"00",
		X"01",X"EF",X"06",X"00",X"EF",X"11",X"00",X"EF",X"13",X"00",X"EF",X"04",X"01",X"EF",X"05",X"01",
		X"EF",X"10",X"13",X"F7",X"43",X"00",X"00",X"21",X"04",X"4E",X"34",X"C9",X"AF",X"32",X"AC",X"4E",
		X"32",X"BC",X"4E",X"3E",X"02",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"3A",X"13",X"4E",X"FE",X"14",
		X"38",X"02",X"3E",X"14",X"E7",X"6F",X"0A",X"08",X"21",X"6F",X"0A",X"6F",X"0A",X"9E",X"21",X"6F",
		X"0A",X"6F",X"0A",X"6F",X"0A",X"97",X"22",X"6F",X"0A",X"6F",X"0A",X"6F",X"0A",X"97",X"22",X"6F",
		X"0A",X"6F",X"0A",X"6F",X"0A",X"97",X"22",X"6F",X"0A",X"6F",X"0A",X"6F",X"0A",X"6F",X"0A",X"21",
		X"04",X"4E",X"34",X"34",X"AF",X"32",X"CC",X"4E",X"32",X"DC",X"4E",X"C9",X"AF",X"32",X"CC",X"4E",
		X"32",X"DC",X"4E",X"06",X"07",X"21",X"0C",X"4E",X"CF",X"CD",X"C9",X"24",X"21",X"04",X"4E",X"34",
		X"21",X"13",X"4E",X"34",X"2A",X"0A",X"4E",X"7E",X"FE",X"14",X"C8",X"23",X"22",X"0A",X"4E",X"C9",
		X"C3",X"88",X"09",X"C3",X"D2",X"09",X"06",X"2E",X"DD",X"21",X"0A",X"4E",X"FD",X"21",X"38",X"4E",
		X"DD",X"56",X"00",X"FD",X"5E",X"00",X"FD",X"72",X"00",X"DD",X"73",X"00",X"DD",X"23",X"FD",X"23",
		X"10",X"EE",X"C9",X"3A",X"A4",X"4D",X"A7",X"C0",X"DD",X"21",X"00",X"4C",X"FD",X"21",X"C8",X"4D",
		X"11",X"00",X"01",X"FD",X"BE",X"00",X"C2",X"D2",X"0B",X"FD",X"36",X"00",X"0E",X"3A",X"A6",X"4D",
		X"A7",X"28",X"1B",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",X"30",X"13",X"21",X"AC",X"4E",X"CB",X"FE",
		X"3E",X"09",X"DD",X"BE",X"0B",X"20",X"04",X"CB",X"BE",X"3E",X"09",X"32",X"0B",X"4C",X"3A",X"A7",
		X"4D",X"A7",X"28",X"1D",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",X"30",X"27",X"3E",X"11",X"DD",X"BE",
		X"03",X"28",X"07",X"DD",X"36",X"03",X"11",X"C3",X"33",X"0B",X"DD",X"36",X"03",X"12",X"C3",X"33",
		X"0B",X"3E",X"01",X"DD",X"BE",X"03",X"28",X"07",X"DD",X"36",X"03",X"01",X"C3",X"33",X"0B",X"DD",
		X"36",X"03",X"01",X"3A",X"A8",X"4D",X"A7",X"28",X"1D",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",X"30",
		X"27",X"3E",X"11",X"DD",X"BE",X"05",X"28",X"07",X"DD",X"36",X"05",X"11",X"C3",X"68",X"0B",X"DD",
		X"36",X"05",X"12",X"C3",X"68",X"0B",X"3E",X"03",X"DD",X"BE",X"05",X"28",X"07",X"DD",X"36",X"05",
		X"03",X"C3",X"68",X"0B",X"DD",X"36",X"05",X"03",X"3A",X"A9",X"4D",X"A7",X"28",X"1D",X"2A",X"CB",
		X"4D",X"A7",X"ED",X"52",X"30",X"27",X"3E",X"11",X"DD",X"BE",X"07",X"28",X"07",X"DD",X"36",X"07",
		X"11",X"C3",X"9D",X"0B",X"DD",X"36",X"07",X"12",X"C3",X"9D",X"0B",X"3E",X"05",X"DD",X"BE",X"07",
		X"28",X"07",X"DD",X"36",X"07",X"05",X"C3",X"9D",X"0B",X"DD",X"36",X"07",X"05",X"3A",X"AA",X"4D",
		X"A7",X"28",X"1D",X"2A",X"CB",X"4D",X"A7",X"ED",X"52",X"30",X"27",X"3E",X"11",X"DD",X"BE",X"09",
		X"28",X"07",X"DD",X"36",X"09",X"11",X"C3",X"D2",X"0B",X"DD",X"36",X"09",X"12",X"C3",X"D2",X"0B",
		X"3E",X"07",X"DD",X"BE",X"09",X"28",X"07",X"DD",X"36",X"09",X"07",X"C3",X"D2",X"0B",X"DD",X"36",
		X"09",X"07",X"FD",X"35",X"00",X"C9",X"06",X"19",X"3A",X"02",X"4E",X"FE",X"22",X"C2",X"E2",X"0B",
		X"06",X"00",X"DD",X"21",X"00",X"4C",X"3A",X"AC",X"4D",X"A7",X"CA",X"F0",X"0B",X"DD",X"70",X"03",
		X"3A",X"AD",X"4D",X"A7",X"CA",X"FA",X"0B",X"DD",X"70",X"05",X"3A",X"AE",X"4D",X"A7",X"CA",X"04",
		X"0C",X"DD",X"70",X"07",X"3A",X"AF",X"4D",X"A7",X"C8",X"DD",X"70",X"09",X"C9",X"21",X"CF",X"4D",
		X"34",X"3E",X"0A",X"BE",X"C0",X"36",X"00",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"15",X"21",X"64",
		X"44",X"3E",X"10",X"BE",X"20",X"02",X"3E",X"00",X"77",X"32",X"78",X"44",X"32",X"84",X"47",X"32",
		X"98",X"47",X"C9",X"21",X"32",X"47",X"3E",X"10",X"BE",X"20",X"02",X"3E",X"00",X"77",X"32",X"78",
		X"46",X"C9",X"3A",X"A4",X"4D",X"A7",X"C0",X"3A",X"94",X"4D",X"07",X"32",X"94",X"4D",X"D0",X"3A",
		X"A0",X"4D",X"A7",X"C2",X"90",X"0C",X"DD",X"21",X"05",X"33",X"FD",X"21",X"00",X"4D",X"CD",X"00",
		X"20",X"22",X"00",X"4D",X"3E",X"03",X"32",X"28",X"4D",X"32",X"2C",X"4D",X"3A",X"00",X"4D",X"FE",
		X"64",X"C2",X"90",X"0C",X"21",X"2C",X"2E",X"22",X"0A",X"4D",X"21",X"00",X"01",X"22",X"14",X"4D",
		X"22",X"1E",X"4D",X"3E",X"02",X"32",X"28",X"4D",X"32",X"2C",X"4D",X"3E",X"01",X"32",X"A0",X"4D",
		X"3A",X"A1",X"4D",X"FE",X"01",X"CA",X"FB",X"0C",X"FE",X"00",X"C2",X"C1",X"0C",X"3A",X"02",X"4D",
		X"FE",X"78",X"CC",X"2E",X"1F",X"FE",X"80",X"CC",X"2E",X"1F",X"3A",X"2D",X"4D",X"32",X"29",X"4D",
		X"DD",X"21",X"20",X"4D",X"FD",X"21",X"02",X"4D",X"CD",X"00",X"20",X"22",X"02",X"4D",X"C3",X"FB",
		X"0C",X"DD",X"21",X"05",X"33",X"FD",X"21",X"02",X"4D",X"CD",X"00",X"20",X"22",X"02",X"4D",X"3E",
		X"03",X"32",X"2D",X"4D",X"32",X"29",X"4D",X"3A",X"02",X"4D",X"FE",X"64",X"C2",X"FB",X"0C",X"21",
		X"2C",X"2E",X"22",X"0C",X"4D",X"21",X"00",X"01",X"22",X"16",X"4D",X"22",X"20",X"4D",X"3E",X"02",
		X"32",X"29",X"4D",X"32",X"2D",X"4D",X"3E",X"01",X"32",X"A1",X"4D",X"3A",X"A2",X"4D",X"FE",X"01",
		X"CA",X"93",X"0D",X"FE",X"00",X"C2",X"2C",X"0D",X"3A",X"04",X"4D",X"FE",X"78",X"CC",X"55",X"1F",
		X"FE",X"80",X"CC",X"55",X"1F",X"3A",X"2E",X"4D",X"32",X"2A",X"4D",X"DD",X"21",X"22",X"4D",X"FD",
		X"21",X"04",X"4D",X"CD",X"00",X"20",X"22",X"04",X"4D",X"C3",X"93",X"0D",X"3A",X"A2",X"4D",X"FE",
		X"03",X"C2",X"59",X"0D",X"DD",X"21",X"FF",X"32",X"FD",X"21",X"04",X"4D",X"CD",X"00",X"20",X"22",
		X"04",X"4D",X"AF",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3A",X"05",X"4D",X"FE",X"80",X"C2",X"93",
		X"0D",X"3E",X"02",X"32",X"A2",X"4D",X"C3",X"93",X"0D",X"DD",X"21",X"05",X"33",X"FD",X"21",X"04",
		X"4D",X"CD",X"00",X"20",X"22",X"04",X"4D",X"3E",X"03",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3A",
		X"04",X"4D",X"FE",X"64",X"C2",X"93",X"0D",X"21",X"2C",X"2E",X"22",X"0E",X"4D",X"21",X"00",X"01",
		X"22",X"18",X"4D",X"22",X"22",X"4D",X"3E",X"02",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"3E",X"01",
		X"32",X"A2",X"4D",X"3A",X"A3",X"4D",X"FE",X"01",X"C8",X"FE",X"00",X"C2",X"C0",X"0D",X"3A",X"06",
		X"4D",X"FE",X"78",X"CC",X"7C",X"1F",X"FE",X"80",X"CC",X"7C",X"1F",X"3A",X"2F",X"4D",X"32",X"2B",
		X"4D",X"DD",X"21",X"24",X"4D",X"FD",X"21",X"06",X"4D",X"CD",X"00",X"20",X"22",X"06",X"4D",X"C9",
		X"3A",X"A3",X"4D",X"FE",X"03",X"C2",X"EA",X"0D",X"DD",X"21",X"03",X"33",X"FD",X"21",X"06",X"4D",
		X"CD",X"00",X"20",X"22",X"06",X"4D",X"3E",X"02",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3A",X"07",
		X"4D",X"FE",X"80",X"C0",X"3E",X"02",X"32",X"A3",X"4D",X"C9",X"DD",X"21",X"05",X"33",X"FD",X"21",
		X"06",X"4D",X"CD",X"00",X"20",X"22",X"06",X"4D",X"3E",X"03",X"32",X"2B",X"4D",X"32",X"2F",X"4D",
		X"3A",X"06",X"4D",X"FE",X"64",X"C0",X"21",X"2C",X"2E",X"22",X"10",X"4D",X"21",X"00",X"01",X"22",
		X"1A",X"4D",X"22",X"24",X"4D",X"3E",X"02",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"3E",X"01",X"32",
		X"A3",X"4D",X"C9",X"21",X"C4",X"4D",X"34",X"3E",X"08",X"BE",X"C0",X"36",X"00",X"3A",X"C0",X"4D",
		X"EE",X"01",X"32",X"C0",X"4D",X"C9",X"3A",X"A6",X"4D",X"A7",X"C0",X"3A",X"C1",X"4D",X"FE",X"07",
		X"C8",X"87",X"2A",X"C2",X"4D",X"23",X"22",X"C2",X"4D",X"5F",X"16",X"00",X"DD",X"21",X"86",X"4D",
		X"DD",X"19",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"A7",X"ED",X"52",X"C0",X"CB",X"3F",X"3C",X"32",
		X"C1",X"4D",X"21",X"01",X"01",X"22",X"B1",X"4D",X"22",X"B3",X"4D",X"C9",X"3A",X"A5",X"4D",X"A7",
		X"28",X"05",X"AF",X"32",X"AC",X"4E",X"C9",X"21",X"AC",X"4E",X"06",X"E0",X"3A",X"0E",X"4E",X"FE",
		X"E4",X"38",X"06",X"78",X"A6",X"CB",X"E7",X"77",X"C9",X"FE",X"D4",X"38",X"06",X"78",X"A6",X"CB",
		X"DF",X"77",X"C9",X"FE",X"B4",X"38",X"06",X"78",X"A6",X"CB",X"D7",X"77",X"C9",X"FE",X"74",X"38",
		X"06",X"78",X"A6",X"CB",X"CF",X"77",X"C9",X"78",X"A6",X"CB",X"C7",X"77",X"C9",X"3A",X"A5",X"4D",
		X"A7",X"C0",X"3A",X"D4",X"4D",X"A7",X"C0",X"3A",X"0E",X"4E",X"FE",X"46",X"28",X"0E",X"FE",X"AA",
		X"C0",X"3A",X"0D",X"4E",X"A7",X"C0",X"21",X"0D",X"4E",X"34",X"18",X"09",X"3A",X"0C",X"4E",X"A7",
		X"C0",X"21",X"0C",X"4E",X"34",X"21",X"94",X"80",X"22",X"D2",X"4D",X"21",X"FD",X"0E",X"3A",X"13",
		X"4E",X"FE",X"14",X"38",X"02",X"3E",X"14",X"47",X"87",X"80",X"D7",X"32",X"0C",X"4C",X"23",X"7E",
		X"32",X"0D",X"4C",X"23",X"7E",X"32",X"D4",X"4D",X"F7",X"8A",X"04",X"00",X"C9",X"00",X"14",X"06",
		X"01",X"0F",X"07",X"02",X"15",X"08",X"02",X"15",X"08",X"04",X"14",X"09",X"04",X"14",X"09",X"05",
		X"17",X"0A",X"05",X"17",X"0A",X"06",X"09",X"0B",X"06",X"09",X"0B",X"03",X"16",X"0C",X"03",X"16",
		X"0C",X"07",X"16",X"0D",X"07",X"16",X"0D",X"07",X"16",X"0D",X"07",X"16",X"0D",X"07",X"16",X"0D",
		X"07",X"16",X"0D",X"07",X"16",X"0D",X"07",X"16",X"0D",X"07",X"16",X"0D",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"36",
		X"AF",X"32",X"D4",X"4D",X"21",X"00",X"00",X"22",X"D2",X"4D",X"C9",X"EF",X"1C",X"9B",X"3A",X"00",
		X"4E",X"3D",X"C8",X"EF",X"1C",X"A2",X"C9",X"CD",X"91",X"12",X"3A",X"A5",X"4D",X"A7",X"C0",X"CD",
		X"66",X"10",X"CD",X"94",X"10",X"CD",X"9E",X"10",X"CD",X"A8",X"10",X"CD",X"B4",X"10",X"3A",X"A4",
		X"4D",X"A7",X"CA",X"39",X"10",X"CD",X"35",X"12",X"C9",X"CD",X"1D",X"17",X"CD",X"89",X"17",X"3A",
		X"A4",X"4D",X"A7",X"C0",X"CD",X"06",X"18",X"CD",X"36",X"1B",X"CD",X"4B",X"1C",X"CD",X"22",X"1D",
		X"CD",X"F9",X"1D",X"3A",X"04",X"4E",X"FE",X"03",X"C0",X"CD",X"76",X"13",X"CD",X"69",X"20",X"CD",
		X"8C",X"20",X"CD",X"AF",X"20",X"C9",X"3A",X"AB",X"4D",X"A7",X"C8",X"3D",X"20",X"08",X"32",X"AB",
		X"4D",X"3C",X"32",X"AC",X"4D",X"C9",X"3D",X"20",X"08",X"32",X"AB",X"4D",X"3C",X"32",X"AD",X"4D",
		X"C9",X"3D",X"20",X"08",X"32",X"AB",X"4D",X"3C",X"32",X"AE",X"4D",X"C9",X"32",X"AF",X"4D",X"3D",
		X"32",X"AB",X"4D",X"C9",X"3A",X"AC",X"4D",X"E7",X"0C",X"00",X"C0",X"10",X"D2",X"10",X"3A",X"AD",
		X"4D",X"E7",X"0C",X"00",X"18",X"11",X"2A",X"11",X"3A",X"AE",X"4D",X"E7",X"0C",X"00",X"5C",X"11",
		X"6E",X"11",X"8F",X"11",X"3A",X"AF",X"4D",X"E7",X"0C",X"00",X"C9",X"11",X"DB",X"11",X"FC",X"11",
		X"CD",X"D8",X"1B",X"2A",X"00",X"4D",X"11",X"64",X"80",X"A7",X"ED",X"52",X"C0",X"21",X"AC",X"4D",
		X"34",X"C9",X"DD",X"21",X"01",X"33",X"FD",X"21",X"00",X"4D",X"CD",X"00",X"20",X"22",X"00",X"4D",
		X"3E",X"01",X"32",X"28",X"4D",X"32",X"2C",X"4D",X"3A",X"00",X"4D",X"FE",X"80",X"C0",X"21",X"2F",
		X"2E",X"22",X"0A",X"4D",X"22",X"31",X"4D",X"AF",X"32",X"A0",X"4D",X"32",X"AC",X"4D",X"32",X"A7",
		X"4D",X"DD",X"21",X"AC",X"4D",X"DD",X"B6",X"00",X"DD",X"B6",X"01",X"DD",X"B6",X"02",X"DD",X"B6",
		X"03",X"C0",X"21",X"AC",X"4E",X"CB",X"B6",X"C9",X"CD",X"AF",X"1C",X"2A",X"02",X"4D",X"11",X"64",
		X"80",X"A7",X"ED",X"52",X"C0",X"21",X"AD",X"4D",X"34",X"C9",X"DD",X"21",X"01",X"33",X"FD",X"21",
		X"02",X"4D",X"CD",X"00",X"20",X"22",X"02",X"4D",X"3E",X"01",X"32",X"29",X"4D",X"32",X"2D",X"4D",
		X"3A",X"02",X"4D",X"FE",X"80",X"C0",X"21",X"2F",X"2E",X"22",X"0C",X"4D",X"22",X"33",X"4D",X"AF",
		X"32",X"A1",X"4D",X"32",X"AD",X"4D",X"32",X"A8",X"4D",X"C3",X"01",X"11",X"CD",X"86",X"1D",X"2A",
		X"04",X"4D",X"11",X"64",X"80",X"A7",X"ED",X"52",X"C0",X"21",X"AE",X"4D",X"34",X"C9",X"DD",X"21",
		X"01",X"33",X"FD",X"21",X"04",X"4D",X"CD",X"00",X"20",X"22",X"04",X"4D",X"3E",X"01",X"32",X"2A",
		X"4D",X"32",X"2E",X"4D",X"3A",X"04",X"4D",X"FE",X"80",X"C0",X"21",X"AE",X"4D",X"34",X"C9",X"DD",
		X"21",X"03",X"33",X"FD",X"21",X"04",X"4D",X"CD",X"00",X"20",X"22",X"04",X"4D",X"3E",X"02",X"32",
		X"2A",X"4D",X"32",X"2E",X"4D",X"3A",X"05",X"4D",X"FE",X"90",X"C0",X"21",X"2F",X"30",X"22",X"0E",
		X"4D",X"22",X"35",X"4D",X"3E",X"01",X"32",X"2A",X"4D",X"32",X"2E",X"4D",X"AF",X"32",X"A2",X"4D",
		X"32",X"AE",X"4D",X"32",X"A9",X"4D",X"C3",X"01",X"11",X"CD",X"5D",X"1E",X"2A",X"06",X"4D",X"11",
		X"64",X"80",X"A7",X"ED",X"52",X"C0",X"21",X"AF",X"4D",X"34",X"C9",X"DD",X"21",X"01",X"33",X"FD",
		X"21",X"06",X"4D",X"CD",X"00",X"20",X"22",X"06",X"4D",X"3E",X"01",X"32",X"2B",X"4D",X"32",X"2F",
		X"4D",X"3A",X"06",X"4D",X"FE",X"80",X"C0",X"21",X"AF",X"4D",X"34",X"C9",X"DD",X"21",X"FF",X"32",
		X"FD",X"21",X"06",X"4D",X"CD",X"00",X"20",X"22",X"06",X"4D",X"AF",X"32",X"2B",X"4D",X"32",X"2F",
		X"4D",X"3A",X"07",X"4D",X"FE",X"70",X"C0",X"21",X"2F",X"2C",X"22",X"10",X"4D",X"22",X"37",X"4D",
		X"3E",X"01",X"32",X"2B",X"4D",X"32",X"2F",X"4D",X"AF",X"32",X"A3",X"4D",X"32",X"AF",X"4D",X"32",
		X"AA",X"4D",X"C3",X"01",X"11",X"3A",X"D1",X"4D",X"E7",X"3F",X"12",X"0C",X"00",X"3F",X"12",X"21",
		X"00",X"4C",X"3A",X"A4",X"4D",X"87",X"5F",X"16",X"00",X"19",X"3A",X"D1",X"4D",X"A7",X"20",X"27",
		X"3A",X"D0",X"4D",X"06",X"27",X"80",X"47",X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"28",
		X"04",X"CB",X"F0",X"CB",X"F8",X"70",X"23",X"36",X"18",X"3E",X"00",X"32",X"0B",X"4C",X"F7",X"4A",
		X"03",X"00",X"21",X"D1",X"4D",X"34",X"C9",X"36",X"20",X"3E",X"09",X"32",X"0B",X"4C",X"3A",X"A4",
		X"4D",X"32",X"AB",X"4D",X"AF",X"32",X"A4",X"4D",X"32",X"D1",X"4D",X"21",X"AC",X"4E",X"CB",X"F6",
		X"C9",X"3A",X"A5",X"4D",X"E7",X"0C",X"00",X"B7",X"12",X"B7",X"12",X"B7",X"12",X"B7",X"12",X"CB",
		X"12",X"F9",X"12",X"06",X"13",X"0E",X"13",X"16",X"13",X"1E",X"13",X"26",X"13",X"2E",X"13",X"36",
		X"13",X"3E",X"13",X"46",X"13",X"53",X"13",X"2A",X"C5",X"4D",X"23",X"22",X"C5",X"4D",X"11",X"78",
		X"00",X"A7",X"ED",X"52",X"C0",X"3E",X"05",X"32",X"A5",X"4D",X"C9",X"21",X"00",X"00",X"CD",X"7E",
		X"26",X"3E",X"34",X"11",X"B4",X"00",X"4F",X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"28",
		X"04",X"3E",X"C0",X"B1",X"4F",X"79",X"32",X"0A",X"4C",X"2A",X"C5",X"4D",X"23",X"22",X"C5",X"4D",
		X"A7",X"ED",X"52",X"C0",X"21",X"A5",X"4D",X"34",X"C9",X"21",X"BC",X"4E",X"CB",X"E6",X"3E",X"35",
		X"11",X"C3",X"00",X"C3",X"D6",X"12",X"3E",X"36",X"11",X"D2",X"00",X"C3",X"D6",X"12",X"3E",X"37",
		X"11",X"E1",X"00",X"C3",X"D6",X"12",X"3E",X"38",X"11",X"F0",X"00",X"C3",X"D6",X"12",X"3E",X"39",
		X"11",X"FF",X"00",X"C3",X"D6",X"12",X"3E",X"3A",X"11",X"0E",X"01",X"C3",X"D6",X"12",X"3E",X"3B",
		X"11",X"1D",X"01",X"C3",X"D6",X"12",X"3E",X"3C",X"11",X"2C",X"01",X"C3",X"D6",X"12",X"3E",X"3D",
		X"11",X"3B",X"01",X"C3",X"D6",X"12",X"21",X"BC",X"4E",X"36",X"20",X"3E",X"3E",X"11",X"59",X"01",
		X"C3",X"D6",X"12",X"3E",X"3F",X"32",X"0A",X"4C",X"2A",X"C5",X"4D",X"23",X"22",X"C5",X"4D",X"11",
		X"B8",X"01",X"A7",X"ED",X"52",X"C0",X"21",X"14",X"4E",X"35",X"21",X"15",X"4E",X"35",X"CD",X"75",
		X"26",X"21",X"04",X"4E",X"34",X"C9",X"3A",X"A6",X"4D",X"A7",X"C8",X"DD",X"21",X"A7",X"4D",X"DD",
		X"7E",X"00",X"DD",X"B6",X"01",X"DD",X"B6",X"02",X"DD",X"B6",X"03",X"CA",X"98",X"13",X"2A",X"CB",
		X"4D",X"2B",X"22",X"CB",X"4D",X"7C",X"B5",X"C0",X"21",X"0B",X"4C",X"36",X"09",X"3A",X"AC",X"4D",
		X"A7",X"C2",X"A7",X"13",X"32",X"A7",X"4D",X"3A",X"AD",X"4D",X"A7",X"C2",X"B1",X"13",X"32",X"A8",
		X"4D",X"3A",X"AE",X"4D",X"A7",X"C2",X"BB",X"13",X"32",X"A9",X"4D",X"3A",X"AF",X"4D",X"A7",X"C2",
		X"C5",X"13",X"32",X"AA",X"4D",X"AF",X"32",X"CB",X"4D",X"32",X"CC",X"4D",X"32",X"A6",X"4D",X"32",
		X"C8",X"4D",X"32",X"D0",X"4D",X"21",X"AC",X"4E",X"CB",X"AE",X"CB",X"BE",X"C9",X"21",X"9E",X"4D",
		X"3A",X"0E",X"4E",X"BE",X"CA",X"EE",X"13",X"21",X"00",X"00",X"22",X"97",X"4D",X"C9",X"2A",X"97",
		X"4D",X"23",X"22",X"97",X"4D",X"ED",X"5B",X"95",X"4D",X"A7",X"ED",X"52",X"C0",X"21",X"00",X"00",
		X"22",X"97",X"4D",X"3A",X"A1",X"4D",X"A7",X"F5",X"CC",X"86",X"20",X"F1",X"C8",X"3A",X"A2",X"4D",
		X"A7",X"F5",X"CC",X"A9",X"20",X"F1",X"C8",X"3A",X"A3",X"4D",X"A7",X"CC",X"D1",X"20",X"C9",X"3A",
		X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"C8",X"47",X"DD",X"21",X"00",X"4C",X"1E",X"08",X"0E",
		X"08",X"16",X"07",X"3A",X"00",X"4D",X"83",X"DD",X"77",X"13",X"3A",X"01",X"4D",X"2F",X"82",X"DD",
		X"77",X"12",X"3A",X"02",X"4D",X"83",X"DD",X"77",X"15",X"3A",X"03",X"4D",X"2F",X"82",X"DD",X"77",
		X"14",X"3A",X"04",X"4D",X"83",X"DD",X"77",X"17",X"3A",X"05",X"4D",X"2F",X"81",X"DD",X"77",X"16",
		X"3A",X"06",X"4D",X"83",X"DD",X"77",X"19",X"3A",X"07",X"4D",X"2F",X"81",X"DD",X"77",X"18",X"3A",
		X"08",X"4D",X"83",X"DD",X"77",X"1B",X"3A",X"09",X"4D",X"2F",X"81",X"DD",X"77",X"1A",X"3A",X"D2",
		X"4D",X"83",X"DD",X"77",X"1D",X"3A",X"D3",X"4D",X"2F",X"81",X"DD",X"77",X"1C",X"C3",X"FE",X"14",
		X"3A",X"72",X"4E",X"47",X"3A",X"09",X"4E",X"A0",X"C0",X"47",X"1E",X"09",X"0E",X"07",X"16",X"06",
		X"DD",X"21",X"00",X"4C",X"3A",X"00",X"4D",X"2F",X"83",X"DD",X"77",X"13",X"3A",X"01",X"4D",X"82",
		X"DD",X"77",X"12",X"3A",X"02",X"4D",X"2F",X"83",X"DD",X"77",X"15",X"3A",X"03",X"4D",X"82",X"DD",
		X"77",X"14",X"3A",X"04",X"4D",X"2F",X"83",X"DD",X"77",X"17",X"3A",X"05",X"4D",X"81",X"DD",X"77",
		X"16",X"3A",X"06",X"4D",X"2F",X"83",X"DD",X"77",X"19",X"3A",X"07",X"4D",X"81",X"DD",X"77",X"18",
		X"3A",X"08",X"4D",X"2F",X"83",X"DD",X"77",X"1B",X"3A",X"09",X"4D",X"81",X"DD",X"77",X"1A",X"3A",
		X"D2",X"4D",X"2F",X"83",X"DD",X"77",X"1D",X"3A",X"D3",X"4D",X"81",X"DD",X"77",X"1C",X"3A",X"A5",
		X"4D",X"A7",X"C2",X"4B",X"15",X"3A",X"A4",X"4D",X"A7",X"C2",X"B4",X"15",X"21",X"1C",X"15",X"E5",
		X"3A",X"30",X"4D",X"E7",X"8C",X"16",X"B1",X"16",X"D6",X"16",X"F7",X"16",X"78",X"A7",X"28",X"2B",
		X"0E",X"C0",X"3A",X"0A",X"4C",X"57",X"A1",X"20",X"05",X"7A",X"B1",X"C3",X"48",X"15",X"3A",X"30",
		X"4D",X"FE",X"02",X"20",X"09",X"CB",X"7A",X"28",X"12",X"7A",X"A9",X"C3",X"48",X"15",X"FE",X"03",
		X"20",X"09",X"CB",X"72",X"28",X"05",X"7A",X"A9",X"32",X"0A",X"4C",X"21",X"C0",X"4D",X"56",X"3E",
		X"1C",X"82",X"DD",X"77",X"02",X"DD",X"77",X"04",X"DD",X"77",X"06",X"DD",X"77",X"08",X"0E",X"20",
		X"3A",X"AC",X"4D",X"A7",X"20",X"06",X"3A",X"A7",X"4D",X"A7",X"20",X"09",X"3A",X"2C",X"4D",X"87",
		X"82",X"81",X"DD",X"77",X"02",X"3A",X"AD",X"4D",X"A7",X"20",X"06",X"3A",X"A8",X"4D",X"A7",X"20",
		X"09",X"3A",X"2D",X"4D",X"87",X"82",X"81",X"DD",X"77",X"04",X"3A",X"AE",X"4D",X"A7",X"20",X"06",
		X"3A",X"A9",X"4D",X"A7",X"20",X"09",X"3A",X"2E",X"4D",X"87",X"82",X"81",X"DD",X"77",X"06",X"3A",
		X"AF",X"4D",X"A7",X"20",X"06",X"3A",X"AA",X"4D",X"A7",X"20",X"09",X"3A",X"2F",X"4D",X"87",X"82",
		X"81",X"DD",X"77",X"08",X"CD",X"E6",X"15",X"CD",X"2D",X"16",X"CD",X"52",X"16",X"78",X"A7",X"C8",
		X"0E",X"C0",X"3A",X"02",X"4C",X"B1",X"32",X"02",X"4C",X"3A",X"04",X"4C",X"B1",X"32",X"04",X"4C",
		X"3A",X"06",X"4C",X"B1",X"32",X"06",X"4C",X"3A",X"08",X"4C",X"B1",X"32",X"08",X"4C",X"3A",X"0C",
		X"4C",X"B1",X"32",X"0C",X"4C",X"C9",X"3A",X"06",X"4E",X"D6",X"05",X"D8",X"3A",X"09",X"4D",X"E6",
		X"0F",X"FE",X"0C",X"38",X"04",X"16",X"18",X"18",X"12",X"FE",X"08",X"38",X"04",X"16",X"14",X"18",
		X"0A",X"FE",X"04",X"38",X"04",X"16",X"10",X"18",X"02",X"16",X"14",X"DD",X"72",X"04",X"14",X"DD",
		X"72",X"06",X"14",X"DD",X"72",X"08",X"14",X"DD",X"72",X"0C",X"DD",X"36",X"0A",X"3F",X"16",X"16",
		X"DD",X"72",X"05",X"DD",X"72",X"07",X"DD",X"72",X"09",X"DD",X"72",X"0D",X"C9",X"3A",X"07",X"4E",
		X"A7",X"C8",X"57",X"3A",X"3A",X"4D",X"D6",X"3D",X"20",X"04",X"DD",X"36",X"0B",X"00",X"7A",X"FE",
		X"0A",X"D8",X"DD",X"36",X"02",X"32",X"DD",X"36",X"03",X"1D",X"FE",X"0C",X"D8",X"DD",X"36",X"02",
		X"33",X"C9",X"3A",X"08",X"4E",X"A7",X"C8",X"57",X"3A",X"3A",X"4D",X"D6",X"3D",X"20",X"04",X"DD",
		X"36",X"0B",X"00",X"7A",X"FE",X"01",X"D8",X"3A",X"C0",X"4D",X"1E",X"08",X"83",X"DD",X"77",X"02",
		X"7A",X"FE",X"03",X"D8",X"3A",X"01",X"4D",X"E6",X"08",X"0F",X"0F",X"0F",X"1E",X"0A",X"83",X"DD",
		X"77",X"0C",X"3C",X"3C",X"DD",X"77",X"02",X"DD",X"36",X"0D",X"1E",X"C9",X"3A",X"09",X"4D",X"E6",
		X"07",X"FE",X"06",X"38",X"05",X"DD",X"36",X"0A",X"30",X"C9",X"FE",X"04",X"38",X"05",X"DD",X"36",
		X"0A",X"2E",X"C9",X"FE",X"02",X"38",X"05",X"DD",X"36",X"0A",X"2C",X"C9",X"DD",X"36",X"0A",X"2E",
		X"C9",X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"06",X"38",X"05",X"DD",X"36",X"0A",X"2F",X"C9",X"FE",
		X"04",X"38",X"05",X"DD",X"36",X"0A",X"2D",X"C9",X"FE",X"02",X"38",X"05",X"DD",X"36",X"0A",X"2F",
		X"C9",X"DD",X"36",X"0A",X"30",X"C9",X"3A",X"09",X"4D",X"E6",X"07",X"FE",X"06",X"38",X"08",X"1E",
		X"2E",X"CB",X"FB",X"DD",X"73",X"0A",X"C9",X"FE",X"04",X"38",X"04",X"1E",X"2C",X"18",X"F2",X"FE",
		X"02",X"30",X"EC",X"1E",X"30",X"18",X"EA",X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"06",X"38",X"05",
		X"DD",X"36",X"0A",X"30",X"C9",X"FE",X"04",X"38",X"08",X"1E",X"2F",X"CB",X"F3",X"DD",X"73",X"0A",
		X"C9",X"FE",X"02",X"38",X"04",X"1E",X"2D",X"18",X"F2",X"1E",X"2F",X"18",X"EE",X"06",X"04",X"ED",
		X"5B",X"39",X"4D",X"3A",X"AF",X"4D",X"A7",X"20",X"09",X"2A",X"37",X"4D",X"A7",X"ED",X"52",X"CA",
		X"63",X"17",X"05",X"3A",X"AE",X"4D",X"A7",X"20",X"09",X"2A",X"35",X"4D",X"A7",X"ED",X"52",X"CA",
		X"63",X"17",X"05",X"3A",X"AD",X"4D",X"A7",X"20",X"09",X"2A",X"33",X"4D",X"A7",X"ED",X"52",X"CA",
		X"63",X"17",X"05",X"3A",X"AC",X"4D",X"A7",X"20",X"09",X"2A",X"31",X"4D",X"A7",X"ED",X"52",X"CA",
		X"63",X"17",X"05",X"78",X"32",X"A4",X"4D",X"32",X"A5",X"4D",X"A7",X"C8",X"21",X"A6",X"4D",X"5F",
		X"16",X"00",X"19",X"7E",X"A7",X"C8",X"AF",X"32",X"A5",X"4D",X"21",X"D0",X"4D",X"34",X"46",X"04",
		X"CD",X"5A",X"2A",X"21",X"BC",X"4E",X"CB",X"DE",X"C9",X"3A",X"A4",X"4D",X"A7",X"C0",X"3A",X"A6",
		X"4D",X"A7",X"C8",X"0E",X"04",X"06",X"04",X"DD",X"21",X"08",X"4D",X"3A",X"AF",X"4D",X"A7",X"20",
		X"13",X"3A",X"06",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"07",X"4D",X"DD",X"96",X"01",
		X"B9",X"DA",X"63",X"17",X"05",X"3A",X"AE",X"4D",X"A7",X"20",X"13",X"3A",X"04",X"4D",X"DD",X"96",
		X"00",X"B9",X"30",X"0A",X"3A",X"05",X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"63",X"17",X"05",X"3A",
		X"AD",X"4D",X"A7",X"20",X"13",X"3A",X"02",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"03",
		X"4D",X"DD",X"96",X"01",X"B9",X"DA",X"63",X"17",X"05",X"3A",X"AC",X"4D",X"A7",X"20",X"13",X"3A",
		X"00",X"4D",X"DD",X"96",X"00",X"B9",X"30",X"0A",X"3A",X"01",X"4D",X"DD",X"96",X"01",X"B9",X"DA",
		X"63",X"17",X"05",X"C3",X"63",X"17",X"21",X"9D",X"4D",X"3E",X"FF",X"BE",X"CA",X"11",X"18",X"35",
		X"C9",X"3A",X"A6",X"4D",X"A7",X"CA",X"2F",X"18",X"2A",X"4C",X"4D",X"29",X"22",X"4C",X"4D",X"2A",
		X"4A",X"4D",X"ED",X"6A",X"22",X"4A",X"4D",X"D0",X"21",X"4C",X"4D",X"34",X"C3",X"43",X"18",X"2A",
		X"48",X"4D",X"29",X"22",X"48",X"4D",X"2A",X"46",X"4D",X"ED",X"6A",X"22",X"46",X"4D",X"D0",X"21",
		X"48",X"4D",X"34",X"3A",X"0E",X"4E",X"32",X"9E",X"4D",X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",
		X"A1",X"4F",X"21",X"3A",X"4D",X"7E",X"06",X"21",X"90",X"38",X"09",X"7E",X"06",X"3B",X"90",X"30",
		X"03",X"C3",X"AB",X"18",X"3E",X"01",X"32",X"BF",X"4D",X"3A",X"00",X"4E",X"FE",X"01",X"CA",X"19",
		X"1A",X"3A",X"04",X"4E",X"FE",X"10",X"D2",X"19",X"1A",X"79",X"A7",X"28",X"06",X"3A",X"40",X"50",
		X"C3",X"86",X"18",X"3A",X"00",X"50",X"CB",X"4F",X"C2",X"99",X"18",X"2A",X"03",X"33",X"3E",X"02",
		X"32",X"30",X"4D",X"22",X"1C",X"4D",X"C3",X"50",X"19",X"CB",X"57",X"C2",X"50",X"19",X"2A",X"FF",
		X"32",X"AF",X"32",X"30",X"4D",X"22",X"1C",X"4D",X"C3",X"50",X"19",X"3A",X"00",X"4E",X"FE",X"01",
		X"CA",X"19",X"1A",X"3A",X"04",X"4E",X"FE",X"10",X"D2",X"19",X"1A",X"79",X"A7",X"28",X"06",X"3A",
		X"40",X"50",X"C3",X"C8",X"18",X"3A",X"00",X"50",X"CB",X"4F",X"CA",X"C9",X"1A",X"CB",X"57",X"CA",
		X"D9",X"1A",X"CB",X"47",X"CA",X"E8",X"1A",X"CB",X"5F",X"CA",X"F8",X"1A",X"2A",X"1C",X"4D",X"22",
		X"26",X"4D",X"06",X"01",X"DD",X"21",X"26",X"4D",X"FD",X"21",X"39",X"4D",X"CD",X"0F",X"20",X"E6",
		X"C0",X"D6",X"C0",X"20",X"4B",X"05",X"C2",X"16",X"19",X"3A",X"30",X"4D",X"0F",X"DA",X"0B",X"19",
		X"3A",X"09",X"4D",X"E6",X"07",X"FE",X"04",X"C8",X"C3",X"40",X"19",X"3A",X"08",X"4D",X"E6",X"07",
		X"FE",X"04",X"C8",X"C3",X"40",X"19",X"DD",X"21",X"1C",X"4D",X"CD",X"0F",X"20",X"E6",X"C0",X"D6",
		X"C0",X"20",X"2D",X"3A",X"30",X"4D",X"0F",X"DA",X"35",X"19",X"3A",X"09",X"4D",X"E6",X"07",X"FE",
		X"04",X"C8",X"C3",X"50",X"19",X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"04",X"C8",X"C3",X"50",X"19",
		X"2A",X"26",X"4D",X"22",X"1C",X"4D",X"05",X"CA",X"50",X"19",X"3A",X"3C",X"4D",X"32",X"30",X"4D",
		X"DD",X"21",X"1C",X"4D",X"FD",X"21",X"08",X"4D",X"CD",X"00",X"20",X"3A",X"30",X"4D",X"0F",X"DA",
		X"75",X"19",X"7D",X"E6",X"07",X"FE",X"04",X"CA",X"85",X"19",X"DA",X"71",X"19",X"2D",X"C3",X"85",
		X"19",X"2C",X"C3",X"85",X"19",X"7C",X"E6",X"07",X"FE",X"04",X"CA",X"85",X"19",X"DA",X"84",X"19",
		X"25",X"C3",X"85",X"19",X"24",X"22",X"08",X"4D",X"CD",X"18",X"20",X"22",X"39",X"4D",X"DD",X"21",
		X"BF",X"4D",X"DD",X"7E",X"00",X"DD",X"36",X"00",X"00",X"A7",X"C0",X"3A",X"D2",X"4D",X"A7",X"28",
		X"2C",X"3A",X"D4",X"4D",X"A7",X"28",X"26",X"2A",X"08",X"4D",X"11",X"94",X"80",X"A7",X"ED",X"52",
		X"20",X"1B",X"06",X"19",X"4F",X"CD",X"42",X"00",X"0E",X"15",X"81",X"4F",X"06",X"1C",X"CD",X"42",
		X"00",X"CD",X"04",X"10",X"F7",X"54",X"05",X"00",X"21",X"BC",X"4E",X"CB",X"D6",X"3E",X"FF",X"32",
		X"9D",X"4D",X"2A",X"39",X"4D",X"CD",X"65",X"00",X"7E",X"FE",X"10",X"28",X"03",X"FE",X"14",X"C0",
		X"DD",X"21",X"0E",X"4E",X"DD",X"34",X"00",X"E6",X"0F",X"CB",X"3F",X"06",X"40",X"70",X"06",X"19",
		X"4F",X"CB",X"39",X"CD",X"42",X"00",X"3C",X"FE",X"01",X"CA",X"FD",X"19",X"87",X"32",X"9D",X"4D",
		X"CD",X"08",X"1B",X"CD",X"6A",X"1A",X"21",X"BC",X"4E",X"3A",X"0E",X"4E",X"0F",X"38",X"05",X"CB",
		X"C6",X"CB",X"8E",X"C9",X"CB",X"86",X"CB",X"CE",X"C9",X"21",X"1C",X"4D",X"7E",X"A7",X"CA",X"2E",
		X"1A",X"3A",X"08",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"38",X"1A",X"C3",X"5C",X"1A",X"3A",X"09",
		X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"5C",X"1A",X"3E",X"05",X"CD",X"D0",X"1E",X"38",X"03",X"EF",
		X"17",X"00",X"DD",X"21",X"26",X"4D",X"FD",X"21",X"12",X"4D",X"CD",X"00",X"20",X"22",X"12",X"4D",
		X"2A",X"26",X"4D",X"22",X"1C",X"4D",X"3A",X"3C",X"4D",X"32",X"30",X"4D",X"DD",X"21",X"1C",X"4D",
		X"FD",X"21",X"08",X"4D",X"CD",X"00",X"20",X"C3",X"85",X"19",X"3A",X"9D",X"4D",X"FE",X"06",X"C0",
		X"2A",X"BD",X"4D",X"22",X"CB",X"4D",X"3E",X"01",X"32",X"A6",X"4D",X"32",X"A7",X"4D",X"32",X"A8",
		X"4D",X"32",X"A9",X"4D",X"32",X"AA",X"4D",X"32",X"B1",X"4D",X"32",X"B2",X"4D",X"32",X"B3",X"4D",
		X"32",X"B4",X"4D",X"32",X"B5",X"4D",X"AF",X"32",X"C8",X"4D",X"32",X"D0",X"4D",X"DD",X"21",X"00",
		X"4C",X"DD",X"36",X"02",X"1C",X"DD",X"36",X"04",X"1C",X"DD",X"36",X"06",X"1C",X"DD",X"36",X"08",
		X"1C",X"DD",X"36",X"03",X"11",X"DD",X"36",X"05",X"11",X"DD",X"36",X"07",X"11",X"DD",X"36",X"09",
		X"11",X"21",X"AC",X"4E",X"CB",X"EE",X"CB",X"BE",X"C9",X"2A",X"03",X"33",X"3E",X"02",X"32",X"3C",
		X"4D",X"22",X"26",X"4D",X"06",X"00",X"C3",X"E4",X"18",X"2A",X"FF",X"32",X"AF",X"32",X"3C",X"4D",
		X"22",X"26",X"4D",X"06",X"00",X"C3",X"E4",X"18",X"2A",X"05",X"33",X"3E",X"03",X"32",X"3C",X"4D",
		X"22",X"26",X"4D",X"06",X"00",X"C3",X"E4",X"18",X"2A",X"01",X"33",X"3E",X"01",X"32",X"3C",X"4D",
		X"22",X"26",X"4D",X"06",X"00",X"C3",X"E4",X"18",X"3A",X"12",X"4E",X"A7",X"CA",X"14",X"1B",X"21",
		X"9F",X"4D",X"34",X"C9",X"3A",X"A3",X"4D",X"A7",X"C0",X"3A",X"A2",X"4D",X"A7",X"CA",X"25",X"1B",
		X"21",X"11",X"4E",X"34",X"C9",X"3A",X"A1",X"4D",X"A7",X"CA",X"31",X"1B",X"21",X"10",X"4E",X"34",
		X"C9",X"21",X"0F",X"4E",X"34",X"C9",X"3A",X"A0",X"4D",X"A7",X"C8",X"3A",X"AC",X"4D",X"A7",X"C0",
		X"CD",X"D7",X"20",X"2A",X"31",X"4D",X"01",X"99",X"4D",X"CD",X"5A",X"20",X"3A",X"99",X"4D",X"A7",
		X"CA",X"6A",X"1B",X"2A",X"60",X"4D",X"29",X"22",X"60",X"4D",X"2A",X"5E",X"4D",X"ED",X"6A",X"22",
		X"5E",X"4D",X"D0",X"21",X"60",X"4D",X"34",X"C3",X"D8",X"1B",X"3A",X"A7",X"4D",X"A7",X"CA",X"88",
		X"1B",X"2A",X"5C",X"4D",X"29",X"22",X"5C",X"4D",X"2A",X"5A",X"4D",X"ED",X"6A",X"22",X"5A",X"4D",
		X"D0",X"21",X"5C",X"4D",X"34",X"C3",X"D8",X"1B",X"3A",X"B7",X"4D",X"A7",X"CA",X"A6",X"1B",X"2A",
		X"50",X"4D",X"29",X"22",X"50",X"4D",X"2A",X"4E",X"4D",X"ED",X"6A",X"22",X"4E",X"4D",X"D0",X"21",
		X"50",X"4D",X"34",X"C3",X"D8",X"1B",X"3A",X"B6",X"4D",X"A7",X"CA",X"C4",X"1B",X"2A",X"54",X"4D",
		X"29",X"22",X"54",X"4D",X"2A",X"52",X"4D",X"ED",X"6A",X"22",X"52",X"4D",X"D0",X"21",X"54",X"4D",
		X"34",X"C3",X"D8",X"1B",X"2A",X"58",X"4D",X"29",X"22",X"58",X"4D",X"2A",X"56",X"4D",X"ED",X"6A",
		X"22",X"56",X"4D",X"D0",X"21",X"58",X"4D",X"34",X"21",X"14",X"4D",X"7E",X"A7",X"CA",X"ED",X"1B",
		X"3A",X"00",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"F7",X"1B",X"C3",X"36",X"1C",X"3A",X"01",X"4D",
		X"E6",X"07",X"FE",X"04",X"C2",X"36",X"1C",X"3E",X"01",X"CD",X"D0",X"1E",X"38",X"1B",X"3A",X"A7",
		X"4D",X"A7",X"CA",X"0B",X"1C",X"EF",X"0C",X"00",X"C3",X"19",X"1C",X"2A",X"0A",X"4D",X"CD",X"52",
		X"20",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"08",X"00",X"CD",X"FE",X"1E",X"DD",X"21",X"1E",X"4D",
		X"FD",X"21",X"0A",X"4D",X"CD",X"00",X"20",X"22",X"0A",X"4D",X"2A",X"1E",X"4D",X"22",X"14",X"4D",
		X"3A",X"2C",X"4D",X"32",X"28",X"4D",X"DD",X"21",X"14",X"4D",X"FD",X"21",X"00",X"4D",X"CD",X"00",
		X"20",X"22",X"00",X"4D",X"CD",X"18",X"20",X"22",X"31",X"4D",X"C9",X"3A",X"A1",X"4D",X"FE",X"01",
		X"C0",X"3A",X"AD",X"4D",X"A7",X"C0",X"2A",X"33",X"4D",X"01",X"9A",X"4D",X"CD",X"5A",X"20",X"3A",
		X"9A",X"4D",X"A7",X"CA",X"7D",X"1C",X"2A",X"6C",X"4D",X"29",X"22",X"6C",X"4D",X"2A",X"6A",X"4D",
		X"ED",X"6A",X"22",X"6A",X"4D",X"D0",X"21",X"6C",X"4D",X"34",X"C3",X"AF",X"1C",X"3A",X"A8",X"4D",
		X"A7",X"CA",X"9B",X"1C",X"2A",X"68",X"4D",X"29",X"22",X"68",X"4D",X"2A",X"66",X"4D",X"ED",X"6A",
		X"22",X"66",X"4D",X"D0",X"21",X"68",X"4D",X"34",X"C3",X"AF",X"1C",X"2A",X"64",X"4D",X"29",X"22",
		X"64",X"4D",X"2A",X"62",X"4D",X"ED",X"6A",X"22",X"62",X"4D",X"D0",X"21",X"64",X"4D",X"34",X"21",
		X"16",X"4D",X"7E",X"A7",X"CA",X"C4",X"1C",X"3A",X"02",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"CE",
		X"1C",X"C3",X"0D",X"1D",X"3A",X"03",X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"0D",X"1D",X"3E",X"02",
		X"CD",X"D0",X"1E",X"38",X"1B",X"3A",X"A8",X"4D",X"A7",X"CA",X"E2",X"1C",X"EF",X"0D",X"00",X"C3",
		X"F0",X"1C",X"2A",X"0C",X"4D",X"CD",X"52",X"20",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"09",X"00",
		X"CD",X"25",X"1F",X"DD",X"21",X"20",X"4D",X"FD",X"21",X"0C",X"4D",X"CD",X"00",X"20",X"22",X"0C",
		X"4D",X"2A",X"20",X"4D",X"22",X"16",X"4D",X"3A",X"2D",X"4D",X"32",X"29",X"4D",X"DD",X"21",X"16",
		X"4D",X"FD",X"21",X"02",X"4D",X"CD",X"00",X"20",X"22",X"02",X"4D",X"CD",X"18",X"20",X"22",X"33",
		X"4D",X"C9",X"3A",X"A2",X"4D",X"FE",X"01",X"C0",X"3A",X"AE",X"4D",X"A7",X"C0",X"2A",X"35",X"4D",
		X"01",X"9B",X"4D",X"CD",X"5A",X"20",X"3A",X"9B",X"4D",X"A7",X"CA",X"54",X"1D",X"2A",X"78",X"4D",
		X"29",X"22",X"78",X"4D",X"2A",X"76",X"4D",X"ED",X"6A",X"22",X"76",X"4D",X"D0",X"21",X"78",X"4D",
		X"34",X"C3",X"86",X"1D",X"3A",X"A9",X"4D",X"A7",X"CA",X"72",X"1D",X"2A",X"74",X"4D",X"29",X"22",
		X"74",X"4D",X"2A",X"72",X"4D",X"ED",X"6A",X"22",X"72",X"4D",X"D0",X"21",X"74",X"4D",X"34",X"C3",
		X"86",X"1D",X"2A",X"70",X"4D",X"29",X"22",X"70",X"4D",X"2A",X"6E",X"4D",X"ED",X"6A",X"22",X"6E",
		X"4D",X"D0",X"21",X"70",X"4D",X"34",X"21",X"18",X"4D",X"7E",X"A7",X"CA",X"9B",X"1D",X"3A",X"04",
		X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"A5",X"1D",X"C3",X"E4",X"1D",X"3A",X"05",X"4D",X"E6",X"07",
		X"FE",X"04",X"C2",X"E4",X"1D",X"3E",X"03",X"CD",X"D0",X"1E",X"38",X"1B",X"3A",X"A9",X"4D",X"A7",
		X"CA",X"B9",X"1D",X"EF",X"0E",X"00",X"C3",X"C7",X"1D",X"2A",X"0E",X"4D",X"CD",X"52",X"20",X"7E",
		X"FE",X"1A",X"28",X"03",X"EF",X"0A",X"00",X"CD",X"4C",X"1F",X"DD",X"21",X"22",X"4D",X"FD",X"21",
		X"0E",X"4D",X"CD",X"00",X"20",X"22",X"0E",X"4D",X"2A",X"22",X"4D",X"22",X"18",X"4D",X"3A",X"2E",
		X"4D",X"32",X"2A",X"4D",X"DD",X"21",X"18",X"4D",X"FD",X"21",X"04",X"4D",X"CD",X"00",X"20",X"22",
		X"04",X"4D",X"CD",X"18",X"20",X"22",X"35",X"4D",X"C9",X"3A",X"A3",X"4D",X"FE",X"01",X"C0",X"3A",
		X"AF",X"4D",X"A7",X"C0",X"2A",X"37",X"4D",X"01",X"9C",X"4D",X"CD",X"5A",X"20",X"3A",X"9C",X"4D",
		X"A7",X"CA",X"2B",X"1E",X"2A",X"84",X"4D",X"29",X"22",X"84",X"4D",X"2A",X"82",X"4D",X"ED",X"6A",
		X"22",X"82",X"4D",X"D0",X"21",X"84",X"4D",X"34",X"C3",X"5D",X"1E",X"3A",X"AA",X"4D",X"A7",X"CA",
		X"49",X"1E",X"2A",X"80",X"4D",X"29",X"22",X"80",X"4D",X"2A",X"7E",X"4D",X"ED",X"6A",X"22",X"7E",
		X"4D",X"D0",X"21",X"80",X"4D",X"34",X"C3",X"5D",X"1E",X"2A",X"7C",X"4D",X"29",X"22",X"7C",X"4D",
		X"2A",X"7A",X"4D",X"ED",X"6A",X"22",X"7A",X"4D",X"D0",X"21",X"7C",X"4D",X"34",X"21",X"1A",X"4D",
		X"7E",X"A7",X"CA",X"72",X"1E",X"3A",X"06",X"4D",X"E6",X"07",X"FE",X"04",X"CA",X"7C",X"1E",X"C3",
		X"BB",X"1E",X"3A",X"07",X"4D",X"E6",X"07",X"FE",X"04",X"C2",X"BB",X"1E",X"3E",X"04",X"CD",X"D0",
		X"1E",X"38",X"1B",X"3A",X"AA",X"4D",X"A7",X"CA",X"90",X"1E",X"EF",X"0F",X"00",X"C3",X"9E",X"1E",
		X"2A",X"10",X"4D",X"CD",X"52",X"20",X"7E",X"FE",X"1A",X"28",X"03",X"EF",X"0B",X"00",X"CD",X"73",
		X"1F",X"DD",X"21",X"24",X"4D",X"FD",X"21",X"10",X"4D",X"CD",X"00",X"20",X"22",X"10",X"4D",X"2A",
		X"24",X"4D",X"22",X"1A",X"4D",X"3A",X"2F",X"4D",X"32",X"2B",X"4D",X"DD",X"21",X"1A",X"4D",X"FD",
		X"21",X"06",X"4D",X"CD",X"00",X"20",X"22",X"06",X"4D",X"CD",X"18",X"20",X"22",X"37",X"4D",X"C9",
		X"87",X"4F",X"06",X"00",X"21",X"09",X"4D",X"09",X"7E",X"FE",X"1D",X"C2",X"E3",X"1E",X"36",X"3D",
		X"C3",X"FC",X"1E",X"FE",X"3E",X"C2",X"ED",X"1E",X"36",X"1E",X"C3",X"FC",X"1E",X"06",X"21",X"90",
		X"DA",X"FC",X"1E",X"7E",X"06",X"3B",X"90",X"D2",X"FC",X"1E",X"A7",X"C9",X"37",X"C9",X"3A",X"B1",
		X"4D",X"A7",X"C8",X"AF",X"32",X"B1",X"4D",X"21",X"FF",X"32",X"3A",X"28",X"4D",X"EE",X"02",X"32",
		X"2C",X"4D",X"47",X"DF",X"22",X"1E",X"4D",X"3A",X"02",X"4E",X"FE",X"22",X"C0",X"22",X"14",X"4D",
		X"78",X"32",X"28",X"4D",X"C9",X"3A",X"B2",X"4D",X"A7",X"C8",X"AF",X"32",X"B2",X"4D",X"21",X"FF",
		X"32",X"3A",X"29",X"4D",X"EE",X"02",X"32",X"2D",X"4D",X"47",X"DF",X"22",X"20",X"4D",X"3A",X"02",
		X"4E",X"FE",X"22",X"C0",X"22",X"16",X"4D",X"78",X"32",X"29",X"4D",X"C9",X"3A",X"B3",X"4D",X"A7",
		X"C8",X"AF",X"32",X"B3",X"4D",X"21",X"FF",X"32",X"3A",X"2A",X"4D",X"EE",X"02",X"32",X"2E",X"4D",
		X"47",X"DF",X"22",X"22",X"4D",X"3A",X"02",X"4E",X"FE",X"22",X"C0",X"22",X"18",X"4D",X"78",X"32",
		X"2A",X"4D",X"C9",X"3A",X"B4",X"4D",X"A7",X"C8",X"AF",X"32",X"B4",X"4D",X"21",X"FF",X"32",X"3A",
		X"2B",X"4D",X"EE",X"02",X"32",X"2F",X"4D",X"47",X"DF",X"22",X"24",X"4D",X"3A",X"02",X"4E",X"FE",
		X"22",X"C0",X"22",X"1A",X"4D",X"78",X"32",X"2B",X"4D",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5D",X"E1",
		X"FD",X"7E",X"00",X"DD",X"86",X"00",X"6F",X"FD",X"7E",X"01",X"DD",X"86",X"01",X"67",X"C9",X"CD",
		X"00",X"20",X"CD",X"65",X"00",X"7E",X"A7",X"C9",X"7D",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",
		X"20",X"6F",X"7C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"1E",X"67",X"C9",X"F5",X"C5",X"7D",
		X"D6",X"20",X"6F",X"7C",X"D6",X"20",X"67",X"06",X"00",X"CB",X"24",X"CB",X"24",X"CB",X"24",X"CB",
		X"24",X"CB",X"10",X"CB",X"24",X"CB",X"10",X"4C",X"26",X"00",X"09",X"01",X"40",X"40",X"09",X"C1",
		X"F1",X"C9",X"CD",X"65",X"00",X"11",X"00",X"04",X"19",X"C9",X"CD",X"52",X"20",X"7E",X"FE",X"1B",
		X"20",X"04",X"3E",X"01",X"02",X"C9",X"AF",X"02",X"C9",X"3A",X"A1",X"4D",X"A7",X"C0",X"3A",X"12",
		X"4E",X"A7",X"CA",X"7E",X"20",X"3A",X"9F",X"4D",X"FE",X"07",X"C0",X"C3",X"86",X"20",X"21",X"B8",
		X"4D",X"3A",X"0F",X"4E",X"BE",X"D8",X"3E",X"02",X"32",X"A1",X"4D",X"C9",X"3A",X"A2",X"4D",X"A7",
		X"C0",X"3A",X"12",X"4E",X"A7",X"CA",X"A1",X"20",X"3A",X"9F",X"4D",X"FE",X"11",X"C0",X"C3",X"A9",
		X"20",X"21",X"B9",X"4D",X"3A",X"10",X"4E",X"BE",X"D8",X"3E",X"03",X"32",X"A2",X"4D",X"C9",X"3A",
		X"A3",X"4D",X"A7",X"C0",X"3A",X"12",X"4E",X"A7",X"CA",X"C9",X"20",X"3A",X"9F",X"4D",X"FE",X"20",
		X"C0",X"AF",X"32",X"12",X"4E",X"32",X"9F",X"4D",X"C9",X"21",X"BA",X"4D",X"3A",X"11",X"4E",X"BE",
		X"D8",X"3E",X"03",X"32",X"A3",X"4D",X"C9",X"3A",X"A3",X"4D",X"A7",X"C8",X"21",X"0E",X"4E",X"3A",
		X"B6",X"4D",X"A7",X"C2",X"F4",X"20",X"3E",X"F4",X"96",X"47",X"3A",X"BB",X"4D",X"90",X"D8",X"3E",
		X"01",X"32",X"B6",X"4D",X"3A",X"B7",X"4D",X"A7",X"C0",X"3E",X"F4",X"96",X"47",X"3A",X"BC",X"4D",
		X"90",X"D8",X"3E",X"01",X"32",X"B7",X"4D",X"C9",X"3A",X"06",X"4E",X"E7",X"1A",X"21",X"40",X"21",
		X"4B",X"21",X"0C",X"00",X"70",X"21",X"7B",X"21",X"86",X"21",X"3A",X"3A",X"4D",X"D6",X"21",X"20",
		X"0F",X"3C",X"32",X"A0",X"4D",X"32",X"B7",X"4D",X"CD",X"06",X"05",X"21",X"06",X"4E",X"34",X"C9",
		X"CD",X"06",X"18",X"CD",X"06",X"18",X"CD",X"36",X"1B",X"CD",X"36",X"1B",X"CD",X"23",X"0E",X"C9",
		X"3A",X"3A",X"4D",X"D6",X"1E",X"C2",X"30",X"21",X"C3",X"2B",X"21",X"3A",X"32",X"4D",X"D6",X"1E",
		X"C2",X"36",X"21",X"CD",X"70",X"1A",X"AF",X"32",X"AC",X"4E",X"32",X"BC",X"4E",X"CD",X"A5",X"05",
		X"22",X"1C",X"4D",X"3A",X"3C",X"4D",X"32",X"30",X"4D",X"F7",X"45",X"07",X"00",X"C3",X"2B",X"21",
		X"3A",X"32",X"4D",X"D6",X"2F",X"C2",X"36",X"21",X"C3",X"2B",X"21",X"3A",X"32",X"4D",X"D6",X"3D",
		X"C2",X"30",X"21",X"C3",X"2B",X"21",X"CD",X"06",X"18",X"CD",X"06",X"18",X"3A",X"3A",X"4D",X"D6",
		X"3D",X"C0",X"32",X"06",X"4E",X"F7",X"45",X"00",X"00",X"21",X"04",X"4E",X"34",X"C9",X"3A",X"07",
		X"4E",X"FD",X"21",X"D2",X"41",X"E7",X"C2",X"21",X"0C",X"00",X"E1",X"21",X"F5",X"21",X"0C",X"22",
		X"1E",X"22",X"44",X"22",X"5D",X"22",X"0C",X"00",X"6A",X"22",X"0C",X"00",X"86",X"22",X"0C",X"00",
		X"8D",X"22",X"3E",X"01",X"32",X"D2",X"45",X"32",X"D3",X"45",X"32",X"F2",X"45",X"32",X"F3",X"45",
		X"CD",X"06",X"05",X"FD",X"36",X"00",X"60",X"FD",X"36",X"01",X"61",X"F7",X"43",X"08",X"00",X"18",
		X"0F",X"3A",X"3A",X"4D",X"D6",X"2C",X"C2",X"30",X"21",X"3C",X"32",X"A0",X"4D",X"32",X"B7",X"4D",
		X"21",X"07",X"4E",X"34",X"C9",X"3A",X"01",X"4D",X"FE",X"77",X"28",X"05",X"FE",X"78",X"C2",X"30",
		X"21",X"21",X"84",X"20",X"22",X"4E",X"4D",X"22",X"50",X"4D",X"18",X"E4",X"3A",X"01",X"4D",X"D6",
		X"78",X"C2",X"37",X"22",X"FD",X"36",X"00",X"62",X"FD",X"36",X"01",X"63",X"18",X"D2",X"3A",X"01",
		X"4D",X"D6",X"7B",X"20",X"12",X"FD",X"36",X"00",X"64",X"FD",X"36",X"01",X"65",X"FD",X"36",X"20",
		X"66",X"FD",X"36",X"21",X"67",X"18",X"B9",X"CD",X"06",X"18",X"CD",X"06",X"18",X"CD",X"36",X"1B",
		X"CD",X"23",X"0E",X"C9",X"3A",X"01",X"4D",X"D6",X"7E",X"20",X"EC",X"FD",X"36",X"00",X"68",X"FD",
		X"36",X"01",X"69",X"FD",X"36",X"20",X"6A",X"FD",X"36",X"21",X"6B",X"18",X"93",X"3A",X"01",X"4D",
		X"D6",X"80",X"20",X"D3",X"F7",X"4F",X"08",X"00",X"18",X"86",X"21",X"01",X"4D",X"34",X"34",X"FD",
		X"36",X"00",X"6C",X"FD",X"36",X"01",X"6D",X"FD",X"36",X"20",X"40",X"FD",X"36",X"21",X"40",X"F7",
		X"4A",X"08",X"00",X"C3",X"F0",X"21",X"F7",X"54",X"08",X"00",X"C3",X"F0",X"21",X"AF",X"32",X"07",
		X"4E",X"21",X"04",X"4E",X"34",X"34",X"C9",X"3A",X"08",X"4E",X"E7",X"A7",X"22",X"BE",X"22",X"0C",
		X"00",X"DD",X"22",X"F5",X"22",X"FE",X"22",X"3A",X"3A",X"4D",X"D6",X"25",X"C2",X"30",X"21",X"3C",
		X"32",X"A0",X"4D",X"32",X"B7",X"4D",X"CD",X"06",X"05",X"21",X"08",X"4E",X"34",X"C9",X"3A",X"01",
		X"4D",X"FE",X"FF",X"28",X"05",X"FE",X"FE",X"C2",X"30",X"21",X"3C",X"3C",X"32",X"01",X"4D",X"3E",
		X"01",X"32",X"B1",X"4D",X"CD",X"FE",X"1E",X"F7",X"4A",X"09",X"00",X"18",X"DC",X"3A",X"32",X"4D",
		X"D6",X"2D",X"28",X"D5",X"3A",X"00",X"4D",X"32",X"D2",X"4D",X"3A",X"01",X"4D",X"D6",X"08",X"32",
		X"D3",X"4D",X"C3",X"30",X"21",X"3A",X"32",X"4D",X"D6",X"1E",X"28",X"BD",X"18",X"E6",X"AF",X"32",
		X"08",X"4E",X"F7",X"45",X"00",X"00",X"21",X"04",X"4E",X"34",X"C9",X"21",X"00",X"50",X"06",X"08",
		X"AF",X"77",X"2C",X"10",X"FC",X"21",X"00",X"40",X"06",X"04",X"32",X"C0",X"50",X"32",X"07",X"50",
		X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F1",X"06",X"04",X"32",X"C0",X"50",X"AF",X"32",
		X"07",X"50",X"3E",X"0F",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F0",X"ED",X"5E",X"3E",X"FA",X"D3",
		X"00",X"AF",X"32",X"07",X"50",X"3C",X"32",X"00",X"50",X"FB",X"76",X"32",X"C0",X"50",X"31",X"C0",
		X"4F",X"AF",X"21",X"00",X"50",X"01",X"08",X"08",X"CF",X"21",X"00",X"4C",X"06",X"BE",X"CF",X"CF",
		X"CF",X"CF",X"21",X"40",X"50",X"06",X"40",X"CF",X"32",X"C0",X"50",X"CD",X"0D",X"24",X"32",X"C0",
		X"50",X"06",X"00",X"CD",X"ED",X"23",X"32",X"C0",X"50",X"21",X"C0",X"4C",X"22",X"80",X"4C",X"22",
		X"82",X"4C",X"3E",X"FF",X"06",X"40",X"CF",X"3E",X"01",X"32",X"00",X"50",X"FB",X"2A",X"82",X"4C",
		X"7E",X"A7",X"FA",X"8D",X"23",X"36",X"FF",X"2C",X"46",X"36",X"FF",X"2C",X"20",X"02",X"2E",X"C0",
		X"22",X"82",X"4C",X"21",X"8D",X"23",X"E5",X"E7",X"ED",X"23",X"D7",X"24",X"19",X"24",X"48",X"24",
		X"3D",X"25",X"8B",X"26",X"0D",X"24",X"98",X"26",X"30",X"27",X"6C",X"27",X"A9",X"27",X"F1",X"27",
		X"3B",X"28",X"65",X"28",X"8F",X"28",X"B9",X"28",X"0D",X"00",X"A2",X"26",X"C9",X"24",X"35",X"2A",
		X"D0",X"26",X"87",X"24",X"E8",X"23",X"E3",X"28",X"E0",X"2A",X"5A",X"2A",X"6A",X"2B",X"EA",X"2B",
		X"5E",X"2C",X"A1",X"2B",X"75",X"26",X"B2",X"26",X"21",X"04",X"4E",X"34",X"C9",X"78",X"E7",X"F3",
		X"23",X"00",X"24",X"3E",X"40",X"01",X"04",X"00",X"21",X"00",X"40",X"CF",X"0D",X"20",X"FC",X"C9",
		X"3E",X"40",X"21",X"40",X"40",X"01",X"04",X"80",X"CF",X"0D",X"20",X"FC",X"C9",X"AF",X"01",X"04",
		X"00",X"21",X"00",X"44",X"CF",X"0D",X"20",X"FC",X"C9",X"21",X"00",X"40",X"01",X"35",X"34",X"0A",
		X"A7",X"C8",X"FA",X"2C",X"24",X"5F",X"16",X"00",X"19",X"2B",X"03",X"0A",X"23",X"77",X"F5",X"E5",
		X"11",X"E0",X"83",X"7D",X"E6",X"1F",X"87",X"26",X"00",X"6F",X"19",X"D1",X"A7",X"ED",X"52",X"F1",
		X"EE",X"01",X"77",X"EB",X"03",X"C3",X"1F",X"24",X"21",X"00",X"40",X"DD",X"21",X"16",X"4E",X"FD",
		X"21",X"B5",X"35",X"16",X"00",X"06",X"1E",X"0E",X"08",X"DD",X"7E",X"00",X"FD",X"5E",X"00",X"19",
		X"07",X"30",X"02",X"36",X"10",X"FD",X"23",X"0D",X"20",X"F2",X"DD",X"23",X"05",X"20",X"E8",X"21",
		X"34",X"4E",X"11",X"64",X"40",X"ED",X"A0",X"11",X"78",X"40",X"ED",X"A0",X"11",X"84",X"43",X"ED",
		X"A0",X"11",X"98",X"43",X"ED",X"A0",X"C9",X"21",X"00",X"40",X"DD",X"21",X"16",X"4E",X"FD",X"21",
		X"B5",X"35",X"16",X"00",X"06",X"1E",X"0E",X"08",X"FD",X"5E",X"00",X"19",X"7E",X"FE",X"10",X"37",
		X"28",X"01",X"3F",X"DD",X"CB",X"00",X"16",X"FD",X"23",X"0D",X"20",X"EC",X"DD",X"23",X"05",X"20",
		X"E5",X"21",X"64",X"40",X"11",X"34",X"4E",X"ED",X"A0",X"21",X"78",X"40",X"ED",X"A0",X"21",X"84",
		X"43",X"ED",X"A0",X"21",X"98",X"43",X"ED",X"A0",X"C9",X"21",X"16",X"4E",X"3E",X"FF",X"06",X"1E",
		X"CF",X"3E",X"14",X"06",X"04",X"CF",X"C9",X"58",X"78",X"FE",X"02",X"3E",X"1F",X"28",X"02",X"3E",
		X"10",X"21",X"40",X"44",X"01",X"04",X"80",X"CF",X"0D",X"20",X"FC",X"3E",X"0F",X"06",X"40",X"21",
		X"C0",X"47",X"CF",X"7B",X"FE",X"01",X"C0",X"3E",X"1A",X"11",X"20",X"00",X"06",X"06",X"DD",X"21",
		X"A0",X"45",X"DD",X"77",X"0C",X"DD",X"77",X"18",X"DD",X"19",X"10",X"F6",X"3E",X"1B",X"06",X"05",
		X"DD",X"21",X"40",X"44",X"DD",X"77",X"0E",X"DD",X"77",X"0F",X"DD",X"77",X"10",X"DD",X"19",X"10",
		X"F3",X"06",X"05",X"DD",X"21",X"20",X"47",X"DD",X"77",X"0E",X"DD",X"77",X"0F",X"DD",X"77",X"10",
		X"DD",X"19",X"10",X"F3",X"3E",X"18",X"32",X"ED",X"45",X"32",X"0D",X"46",X"C9",X"DD",X"21",X"00",
		X"4C",X"DD",X"36",X"02",X"20",X"DD",X"36",X"04",X"20",X"DD",X"36",X"06",X"20",X"DD",X"36",X"08",
		X"20",X"DD",X"36",X"0A",X"2C",X"DD",X"36",X"0C",X"3F",X"DD",X"36",X"03",X"01",X"DD",X"36",X"05",
		X"03",X"DD",X"36",X"07",X"05",X"DD",X"36",X"09",X"07",X"DD",X"36",X"0B",X"09",X"DD",X"36",X"0D",
		X"00",X"78",X"A7",X"C2",X"0F",X"26",X"21",X"64",X"80",X"22",X"00",X"4D",X"21",X"7C",X"80",X"22",
		X"02",X"4D",X"21",X"7C",X"90",X"22",X"04",X"4D",X"21",X"7C",X"70",X"22",X"06",X"4D",X"21",X"C4",
		X"80",X"22",X"08",X"4D",X"21",X"2C",X"2E",X"22",X"0A",X"4D",X"22",X"31",X"4D",X"21",X"2F",X"2E",
		X"22",X"0C",X"4D",X"22",X"33",X"4D",X"21",X"2F",X"30",X"22",X"0E",X"4D",X"22",X"35",X"4D",X"21",
		X"2F",X"2C",X"22",X"10",X"4D",X"22",X"37",X"4D",X"21",X"38",X"2E",X"22",X"12",X"4D",X"22",X"39",
		X"4D",X"21",X"00",X"01",X"22",X"14",X"4D",X"22",X"1E",X"4D",X"21",X"01",X"00",X"22",X"16",X"4D",
		X"22",X"20",X"4D",X"21",X"FF",X"00",X"22",X"18",X"4D",X"22",X"22",X"4D",X"21",X"FF",X"00",X"22",
		X"1A",X"4D",X"22",X"24",X"4D",X"21",X"00",X"01",X"22",X"1C",X"4D",X"22",X"26",X"4D",X"21",X"02",
		X"01",X"22",X"28",X"4D",X"22",X"2C",X"4D",X"21",X"03",X"03",X"22",X"2A",X"4D",X"22",X"2E",X"4D",
		X"3E",X"02",X"32",X"30",X"4D",X"32",X"3C",X"4D",X"21",X"00",X"00",X"22",X"D2",X"4D",X"C9",X"21",
		X"94",X"00",X"22",X"00",X"4D",X"22",X"02",X"4D",X"22",X"04",X"4D",X"22",X"06",X"4D",X"21",X"32",
		X"1E",X"22",X"0A",X"4D",X"22",X"0C",X"4D",X"22",X"0E",X"4D",X"22",X"10",X"4D",X"22",X"31",X"4D",
		X"22",X"33",X"4D",X"22",X"35",X"4D",X"22",X"37",X"4D",X"21",X"00",X"01",X"22",X"14",X"4D",X"22",
		X"16",X"4D",X"22",X"18",X"4D",X"22",X"1A",X"4D",X"22",X"1E",X"4D",X"22",X"20",X"4D",X"22",X"22",
		X"4D",X"22",X"24",X"4D",X"22",X"1C",X"4D",X"22",X"26",X"4D",X"21",X"28",X"4D",X"3E",X"02",X"06",
		X"09",X"CF",X"32",X"3C",X"4D",X"21",X"94",X"08",X"22",X"08",X"4D",X"21",X"32",X"1F",X"22",X"12",
		X"4D",X"22",X"39",X"4D",X"C9",X"21",X"00",X"00",X"22",X"D2",X"4D",X"22",X"08",X"4D",X"22",X"00",
		X"4D",X"22",X"02",X"4D",X"22",X"04",X"4D",X"22",X"06",X"4D",X"C9",X"3E",X"55",X"32",X"94",X"4D",
		X"05",X"C8",X"3E",X"01",X"32",X"A0",X"4D",X"C9",X"3E",X"01",X"32",X"00",X"4E",X"AF",X"32",X"01",
		X"4E",X"C9",X"AF",X"11",X"00",X"4D",X"21",X"00",X"4E",X"12",X"13",X"A7",X"ED",X"52",X"C2",X"A6",
		X"26",X"C9",X"DD",X"21",X"36",X"41",X"3A",X"71",X"4E",X"E6",X"0F",X"C6",X"30",X"DD",X"77",X"00",
		X"3A",X"71",X"4E",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"C8",X"C6",X"30",X"DD",X"77",X"20",X"C9",
		X"3A",X"80",X"50",X"47",X"E6",X"03",X"C2",X"DE",X"26",X"21",X"6E",X"4E",X"36",X"FF",X"4F",X"1F",
		X"CE",X"00",X"32",X"6B",X"4E",X"E6",X"02",X"A9",X"32",X"6D",X"4E",X"78",X"0F",X"0F",X"E6",X"03",
		X"3C",X"FE",X"04",X"20",X"01",X"3C",X"32",X"6F",X"4E",X"78",X"0F",X"0F",X"0F",X"0F",X"E6",X"03",
		X"21",X"28",X"27",X"D7",X"32",X"71",X"4E",X"78",X"07",X"2F",X"E6",X"01",X"32",X"75",X"4E",X"78",
		X"07",X"07",X"2F",X"E6",X"01",X"47",X"21",X"2C",X"27",X"DF",X"22",X"73",X"4E",X"3A",X"40",X"50",
		X"07",X"2F",X"E6",X"01",X"32",X"72",X"4E",X"C9",X"10",X"15",X"20",X"FF",X"68",X"00",X"7D",X"00",
		X"3A",X"C1",X"4D",X"CB",X"47",X"C2",X"58",X"27",X"3A",X"B6",X"4D",X"A7",X"20",X"1A",X"3A",X"04",
		X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0A",X"4D",X"3A",X"2C",X"4D",X"11",X"1D",X"22",X"CD",X"66",
		X"29",X"22",X"1E",X"4D",X"32",X"2C",X"4D",X"C9",X"2A",X"0A",X"4D",X"ED",X"5B",X"39",X"4D",X"3A",
		X"2C",X"4D",X"CD",X"66",X"29",X"22",X"1E",X"4D",X"32",X"2C",X"4D",X"C9",X"3A",X"C1",X"4D",X"CB",
		X"47",X"C2",X"8E",X"27",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0C",X"4D",X"3A",X"2D",
		X"4D",X"11",X"1D",X"39",X"CD",X"66",X"29",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"ED",X"5B",
		X"39",X"4D",X"2A",X"1C",X"4D",X"29",X"29",X"19",X"EB",X"2A",X"0C",X"4D",X"3A",X"2D",X"4D",X"CD",
		X"66",X"29",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"3A",X"C1",X"4D",X"CB",X"47",X"C2",X"CB",
		X"27",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",X"11",X"40",
		X"20",X"CD",X"66",X"29",X"22",X"22",X"4D",X"32",X"2E",X"4D",X"C9",X"ED",X"4B",X"0A",X"4D",X"ED",
		X"5B",X"39",X"4D",X"2A",X"1C",X"4D",X"29",X"19",X"7D",X"87",X"91",X"6F",X"7C",X"87",X"90",X"67",
		X"EB",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",X"CD",X"66",X"29",X"22",X"22",X"4D",X"32",X"2E",X"4D",
		X"C9",X"3A",X"C1",X"4D",X"CB",X"47",X"C2",X"13",X"28",X"3A",X"04",X"4E",X"FE",X"03",X"20",X"13",
		X"2A",X"10",X"4D",X"3A",X"2F",X"4D",X"11",X"40",X"3B",X"CD",X"66",X"29",X"22",X"24",X"4D",X"32",
		X"2F",X"4D",X"C9",X"DD",X"21",X"39",X"4D",X"FD",X"21",X"10",X"4D",X"CD",X"EA",X"29",X"11",X"40",
		X"00",X"A7",X"ED",X"52",X"DA",X"00",X"28",X"2A",X"10",X"4D",X"ED",X"5B",X"39",X"4D",X"3A",X"2F",
		X"4D",X"CD",X"66",X"29",X"22",X"24",X"4D",X"32",X"2F",X"4D",X"C9",X"3A",X"AC",X"4D",X"A7",X"CA",
		X"55",X"28",X"11",X"2C",X"2E",X"2A",X"0A",X"4D",X"3A",X"2C",X"4D",X"CD",X"66",X"29",X"22",X"1E",
		X"4D",X"32",X"2C",X"4D",X"C9",X"2A",X"0A",X"4D",X"3A",X"2C",X"4D",X"CD",X"1E",X"29",X"22",X"1E",
		X"4D",X"32",X"2C",X"4D",X"C9",X"3A",X"AD",X"4D",X"A7",X"CA",X"7F",X"28",X"11",X"2C",X"2E",X"2A",
		X"0C",X"4D",X"3A",X"2D",X"4D",X"CD",X"66",X"29",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"2A",
		X"0C",X"4D",X"3A",X"2D",X"4D",X"CD",X"1E",X"29",X"22",X"20",X"4D",X"32",X"2D",X"4D",X"C9",X"3A",
		X"AE",X"4D",X"A7",X"CA",X"A9",X"28",X"11",X"2C",X"2E",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",X"CD",
		X"66",X"29",X"22",X"22",X"4D",X"32",X"2E",X"4D",X"C9",X"2A",X"0E",X"4D",X"3A",X"2E",X"4D",X"CD",
		X"1E",X"29",X"22",X"22",X"4D",X"32",X"2E",X"4D",X"C9",X"3A",X"AF",X"4D",X"A7",X"CA",X"D3",X"28",
		X"11",X"2C",X"2E",X"2A",X"10",X"4D",X"3A",X"2F",X"4D",X"CD",X"66",X"29",X"22",X"24",X"4D",X"32",
		X"2F",X"4D",X"C9",X"2A",X"10",X"4D",X"3A",X"2F",X"4D",X"CD",X"1E",X"29",X"22",X"24",X"4D",X"32",
		X"2F",X"4D",X"C9",X"3A",X"A7",X"4D",X"A7",X"CA",X"FE",X"28",X"2A",X"12",X"4D",X"ED",X"5B",X"0C",
		X"4D",X"3A",X"3C",X"4D",X"CD",X"66",X"29",X"22",X"26",X"4D",X"32",X"3C",X"4D",X"C9",X"2A",X"39",
		X"4D",X"ED",X"4B",X"0C",X"4D",X"7D",X"87",X"91",X"6F",X"7C",X"87",X"90",X"67",X"EB",X"2A",X"12",
		X"4D",X"3A",X"3C",X"4D",X"CD",X"66",X"29",X"22",X"26",X"4D",X"32",X"3C",X"4D",X"C9",X"22",X"3E",
		X"4D",X"EE",X"02",X"32",X"3D",X"4D",X"CD",X"23",X"2A",X"E6",X"03",X"21",X"3B",X"4D",X"77",X"87",
		X"5F",X"16",X"00",X"DD",X"21",X"FF",X"32",X"DD",X"19",X"FD",X"21",X"3E",X"4D",X"3A",X"3D",X"4D",
		X"BE",X"CA",X"57",X"29",X"CD",X"0F",X"20",X"E6",X"C0",X"D6",X"C0",X"28",X"0A",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"3A",X"3B",X"4D",X"C9",X"DD",X"23",X"DD",X"23",X"21",X"3B",X"4D",X"7E",X"3C",
		X"E6",X"03",X"77",X"C3",X"3D",X"29",X"22",X"3E",X"4D",X"ED",X"53",X"40",X"4D",X"32",X"3B",X"4D",
		X"EE",X"02",X"32",X"3D",X"4D",X"21",X"FF",X"FF",X"22",X"44",X"4D",X"DD",X"21",X"FF",X"32",X"FD",
		X"21",X"3E",X"4D",X"21",X"C7",X"4D",X"36",X"00",X"3A",X"3D",X"4D",X"BE",X"CA",X"C6",X"29",X"CD",
		X"00",X"20",X"22",X"42",X"4D",X"CD",X"65",X"00",X"7E",X"E6",X"C0",X"D6",X"C0",X"28",X"27",X"DD",
		X"E5",X"FD",X"E5",X"DD",X"21",X"40",X"4D",X"FD",X"21",X"42",X"4D",X"CD",X"EA",X"29",X"FD",X"E1",
		X"DD",X"E1",X"EB",X"2A",X"44",X"4D",X"A7",X"ED",X"52",X"DA",X"C6",X"29",X"ED",X"53",X"44",X"4D",
		X"3A",X"C7",X"4D",X"32",X"3B",X"4D",X"DD",X"23",X"DD",X"23",X"21",X"C7",X"4D",X"34",X"3E",X"04",
		X"BE",X"C2",X"88",X"29",X"3A",X"3B",X"4D",X"87",X"5F",X"16",X"00",X"DD",X"21",X"FF",X"32",X"DD",
		X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"CB",X"3F",X"C9",X"DD",X"7E",X"00",X"FD",X"46",X"00",
		X"90",X"D2",X"F9",X"29",X"78",X"DD",X"46",X"00",X"90",X"CD",X"12",X"2A",X"E5",X"DD",X"7E",X"01",
		X"FD",X"46",X"01",X"90",X"D2",X"0C",X"2A",X"78",X"DD",X"46",X"01",X"90",X"CD",X"12",X"2A",X"C1",
		X"09",X"C9",X"67",X"5F",X"2E",X"00",X"55",X"0E",X"08",X"29",X"D2",X"1E",X"2A",X"19",X"0D",X"C2",
		X"19",X"2A",X"C9",X"2A",X"C9",X"4D",X"54",X"5D",X"29",X"29",X"19",X"23",X"7C",X"E6",X"1F",X"67",
		X"7E",X"22",X"C9",X"4D",X"C9",X"11",X"40",X"40",X"21",X"C0",X"43",X"A7",X"ED",X"52",X"C8",X"1A",
		X"FE",X"10",X"CA",X"53",X"2A",X"FE",X"12",X"CA",X"53",X"2A",X"FE",X"14",X"CA",X"53",X"2A",X"13",
		X"C3",X"38",X"2A",X"3E",X"40",X"12",X"13",X"C3",X"38",X"2A",X"3A",X"00",X"4E",X"FE",X"01",X"C8",
		X"21",X"17",X"2B",X"DF",X"EB",X"CD",X"0B",X"2B",X"7B",X"86",X"27",X"77",X"23",X"7A",X"8E",X"27",
		X"77",X"5F",X"23",X"3E",X"00",X"8E",X"27",X"77",X"57",X"EB",X"29",X"29",X"29",X"29",X"3A",X"71",
		X"4E",X"3D",X"BC",X"DC",X"33",X"2B",X"CD",X"AF",X"2A",X"13",X"13",X"13",X"21",X"8A",X"4E",X"06",
		X"03",X"1A",X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"CD",X"0B",X"2B",X"11",X"88",
		X"4E",X"01",X"03",X"00",X"ED",X"B0",X"1B",X"01",X"04",X"03",X"21",X"F2",X"43",X"18",X"0F",X"3A",
		X"09",X"4E",X"01",X"04",X"03",X"21",X"FC",X"43",X"A7",X"28",X"03",X"21",X"E9",X"43",X"1A",X"0F",
		X"0F",X"0F",X"0F",X"CD",X"CE",X"2A",X"1A",X"CD",X"CE",X"2A",X"1B",X"10",X"F1",X"C9",X"E6",X"0F",
		X"28",X"04",X"0E",X"00",X"18",X"07",X"79",X"A7",X"28",X"03",X"3E",X"40",X"0D",X"77",X"2B",X"C9",
		X"06",X"00",X"CD",X"5E",X"2C",X"AF",X"21",X"80",X"4E",X"06",X"08",X"CF",X"01",X"04",X"03",X"11",
		X"82",X"4E",X"21",X"FC",X"43",X"CD",X"BE",X"2A",X"01",X"04",X"03",X"11",X"86",X"4E",X"21",X"E9",
		X"43",X"3A",X"70",X"4E",X"A7",X"20",X"B7",X"0E",X"06",X"18",X"B3",X"3A",X"09",X"4E",X"21",X"80",
		X"4E",X"A7",X"C8",X"21",X"84",X"4E",X"C9",X"10",X"00",X"50",X"00",X"00",X"02",X"00",X"04",X"00",
		X"08",X"00",X"16",X"00",X"01",X"00",X"03",X"00",X"05",X"00",X"07",X"00",X"10",X"00",X"20",X"00",
		X"30",X"00",X"50",X"13",X"6B",X"62",X"1B",X"CB",X"46",X"C0",X"CB",X"C6",X"21",X"9C",X"4E",X"CB",
		X"C6",X"21",X"14",X"4E",X"34",X"21",X"15",X"4E",X"34",X"46",X"21",X"1A",X"40",X"0E",X"05",X"78",
		X"A7",X"28",X"0E",X"FE",X"06",X"30",X"0A",X"3E",X"20",X"CD",X"8F",X"2B",X"2B",X"2B",X"0D",X"10",
		X"F6",X"0D",X"F8",X"CD",X"7E",X"2B",X"2B",X"2B",X"18",X"F7",X"3A",X"00",X"4E",X"FE",X"01",X"C8",
		X"CD",X"CD",X"2B",X"12",X"44",X"09",X"0A",X"02",X"21",X"15",X"4E",X"46",X"18",X"CC",X"3E",X"40",
		X"E5",X"D5",X"77",X"23",X"77",X"11",X"1F",X"00",X"19",X"77",X"23",X"77",X"D1",X"E1",X"C9",X"E5",
		X"D5",X"11",X"1F",X"00",X"77",X"3C",X"23",X"77",X"3C",X"19",X"77",X"3C",X"23",X"77",X"D1",X"E1",
		X"C9",X"3A",X"6E",X"4E",X"FE",X"FF",X"20",X"05",X"06",X"02",X"C3",X"5E",X"2C",X"06",X"01",X"CD",
		X"5E",X"2C",X"3A",X"6E",X"4E",X"E6",X"F0",X"28",X"09",X"0F",X"0F",X"0F",X"0F",X"C6",X"30",X"32",
		X"34",X"40",X"3A",X"6E",X"4E",X"E6",X"0F",X"C6",X"30",X"32",X"33",X"40",X"C9",X"E1",X"5E",X"23",
		X"56",X"23",X"4E",X"23",X"46",X"23",X"7E",X"23",X"E5",X"EB",X"11",X"20",X"00",X"E5",X"C5",X"71",
		X"23",X"10",X"FC",X"C1",X"E1",X"19",X"3D",X"20",X"F4",X"C9",X"3A",X"00",X"4E",X"FE",X"01",X"C8",
		X"3A",X"13",X"4E",X"3C",X"FE",X"08",X"D2",X"2E",X"2C",X"11",X"08",X"3B",X"47",X"0E",X"07",X"21",
		X"04",X"40",X"1A",X"CD",X"8F",X"2B",X"3E",X"04",X"84",X"67",X"13",X"1A",X"CD",X"80",X"2B",X"3E",
		X"FC",X"84",X"67",X"13",X"23",X"23",X"0D",X"10",X"E9",X"0D",X"F8",X"CD",X"7E",X"2B",X"3E",X"04",
		X"84",X"67",X"AF",X"CD",X"80",X"2B",X"3E",X"FC",X"84",X"67",X"23",X"23",X"18",X"EB",X"FE",X"13",
		X"38",X"02",X"3E",X"13",X"D6",X"07",X"4F",X"06",X"00",X"21",X"08",X"3B",X"09",X"09",X"EB",X"06",
		X"07",X"C3",X"FD",X"2B",X"47",X"E6",X"0F",X"C6",X"00",X"27",X"4F",X"78",X"E6",X"F0",X"28",X"0B",
		X"0F",X"0F",X"0F",X"0F",X"47",X"AF",X"C6",X"16",X"27",X"10",X"FB",X"81",X"27",X"C9",X"21",X"A5",
		X"36",X"DF",X"5E",X"23",X"56",X"DD",X"21",X"00",X"44",X"DD",X"19",X"DD",X"E5",X"11",X"00",X"FC",
		X"DD",X"19",X"11",X"FF",X"FF",X"CB",X"7E",X"20",X"03",X"11",X"E0",X"FF",X"23",X"78",X"01",X"00",
		X"00",X"87",X"38",X"28",X"7E",X"FE",X"2F",X"28",X"09",X"DD",X"77",X"00",X"23",X"DD",X"19",X"04",
		X"18",X"F2",X"23",X"DD",X"E1",X"7E",X"A7",X"FA",X"A4",X"2C",X"7E",X"DD",X"77",X"00",X"23",X"DD",
		X"19",X"10",X"F7",X"C9",X"DD",X"77",X"00",X"DD",X"19",X"10",X"F9",X"C9",X"7E",X"FE",X"2F",X"28",
		X"0A",X"DD",X"36",X"00",X"40",X"23",X"DD",X"19",X"04",X"18",X"F1",X"23",X"04",X"ED",X"B1",X"18",
		X"D2",X"21",X"C8",X"3B",X"DD",X"21",X"CC",X"4E",X"FD",X"21",X"8C",X"4E",X"CD",X"44",X"2D",X"47",
		X"3A",X"CC",X"4E",X"A7",X"28",X"04",X"78",X"32",X"91",X"4E",X"21",X"CC",X"3B",X"DD",X"21",X"DC",
		X"4E",X"FD",X"21",X"92",X"4E",X"CD",X"44",X"2D",X"47",X"3A",X"DC",X"4E",X"A7",X"28",X"04",X"78",
		X"32",X"96",X"4E",X"21",X"D0",X"3B",X"DD",X"21",X"EC",X"4E",X"FD",X"21",X"97",X"4E",X"CD",X"44",
		X"2D",X"47",X"3A",X"EC",X"4E",X"A7",X"C8",X"78",X"32",X"9B",X"4E",X"C9",X"21",X"30",X"3B",X"DD",
		X"21",X"9C",X"4E",X"FD",X"21",X"8C",X"4E",X"CD",X"EE",X"2D",X"32",X"91",X"4E",X"21",X"40",X"3B",
		X"DD",X"21",X"AC",X"4E",X"FD",X"21",X"92",X"4E",X"CD",X"EE",X"2D",X"32",X"96",X"4E",X"21",X"80",
		X"3B",X"DD",X"21",X"BC",X"4E",X"FD",X"21",X"97",X"4E",X"CD",X"EE",X"2D",X"32",X"9B",X"4E",X"AF",
		X"32",X"90",X"4E",X"C9",X"DD",X"7E",X"00",X"A7",X"CA",X"F4",X"2D",X"4F",X"06",X"08",X"1E",X"80",
		X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",X"DD",X"7E",X"02",X"A3",X"20",X"07",X"DD",
		X"73",X"02",X"05",X"DF",X"18",X"0C",X"DD",X"35",X"0C",X"C2",X"D7",X"2D",X"DD",X"6E",X"06",X"DD",
		X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"FE",X"F0",X"38",X"27",X"21",X"6C",
		X"2D",X"E5",X"E6",X"0F",X"E7",X"55",X"2F",X"65",X"2F",X"77",X"2F",X"89",X"2F",X"9B",X"2F",X"0C",
		X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",X"00",X"0C",
		X"00",X"0C",X"00",X"AD",X"2F",X"47",X"E6",X"1F",X"28",X"03",X"DD",X"70",X"0D",X"DD",X"4E",X"09",
		X"DD",X"7E",X"0B",X"E6",X"08",X"28",X"02",X"0E",X"00",X"DD",X"71",X"0F",X"78",X"07",X"07",X"07",
		X"E6",X"07",X"21",X"B0",X"3B",X"D7",X"DD",X"77",X"0C",X"78",X"E6",X"1F",X"28",X"09",X"E6",X"0F",
		X"21",X"B8",X"3B",X"D7",X"DD",X"77",X"0E",X"DD",X"6E",X"0E",X"26",X"00",X"DD",X"7E",X"0D",X"E6",
		X"10",X"28",X"02",X"3E",X"01",X"DD",X"86",X"04",X"CA",X"E8",X"2E",X"C3",X"E4",X"2E",X"DD",X"7E",
		X"00",X"A7",X"20",X"27",X"DD",X"7E",X"02",X"A7",X"C8",X"DD",X"36",X"02",X"00",X"DD",X"36",X"0D",
		X"00",X"DD",X"36",X"0E",X"00",X"DD",X"36",X"0F",X"00",X"FD",X"36",X"00",X"00",X"FD",X"36",X"01",
		X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",X"00",X"AF",X"C9",X"4F",X"06",X"08",X"1E",X"80",
		X"7B",X"A1",X"20",X"05",X"CB",X"3B",X"10",X"F8",X"C9",X"DD",X"7E",X"02",X"A3",X"20",X"3F",X"DD",
		X"73",X"02",X"05",X"78",X"07",X"07",X"07",X"4F",X"06",X"00",X"E5",X"09",X"DD",X"E5",X"D1",X"13",
		X"13",X"13",X"01",X"08",X"00",X"ED",X"B0",X"E1",X"DD",X"7E",X"06",X"E6",X"7F",X"DD",X"77",X"0C",
		X"DD",X"7E",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",X"47",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",
		X"DD",X"77",X"0B",X"E6",X"08",X"20",X"07",X"DD",X"70",X"0F",X"DD",X"36",X"0D",X"00",X"DD",X"35",
		X"0C",X"20",X"5A",X"DD",X"7E",X"08",X"A7",X"28",X"10",X"DD",X"35",X"08",X"20",X"0B",X"7B",X"2F",
		X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"EE",X"2D",X"DD",X"7E",X"06",X"E6",X"7F",X"DD",X"77",
		X"0C",X"DD",X"CB",X"06",X"7E",X"28",X"16",X"DD",X"7E",X"05",X"ED",X"44",X"DD",X"77",X"05",X"DD",
		X"CB",X"0D",X"46",X"DD",X"CB",X"0D",X"C6",X"28",X"24",X"DD",X"CB",X"0D",X"86",X"DD",X"7E",X"04",
		X"DD",X"86",X"07",X"DD",X"77",X"04",X"DD",X"77",X"0E",X"DD",X"7E",X"09",X"DD",X"86",X"0A",X"DD",
		X"77",X"09",X"47",X"DD",X"7E",X"0B",X"E6",X"08",X"20",X"03",X"DD",X"70",X"0F",X"DD",X"7E",X"0E",
		X"DD",X"86",X"05",X"DD",X"77",X"0E",X"6F",X"26",X"00",X"DD",X"7E",X"03",X"E6",X"70",X"28",X"08",
		X"0F",X"0F",X"0F",X"0F",X"47",X"29",X"10",X"FD",X"FD",X"75",X"00",X"7D",X"0F",X"0F",X"0F",X"0F",
		X"FD",X"77",X"01",X"FD",X"74",X"02",X"7C",X"0F",X"0F",X"0F",X"0F",X"FD",X"77",X"03",X"DD",X"7E",
		X"0B",X"E7",X"22",X"2F",X"26",X"2F",X"2B",X"2F",X"3C",X"2F",X"43",X"2F",X"4A",X"2F",X"4B",X"2F",
		X"4C",X"2F",X"4D",X"2F",X"4E",X"2F",X"4F",X"2F",X"50",X"2F",X"51",X"2F",X"52",X"2F",X"53",X"2F",
		X"54",X"2F",X"DD",X"7E",X"0F",X"C9",X"DD",X"7E",X"0F",X"18",X"09",X"3A",X"84",X"4C",X"E6",X"01",
		X"DD",X"7E",X"0F",X"C0",X"E6",X"0F",X"C8",X"3D",X"DD",X"77",X"0F",X"C9",X"3A",X"84",X"4C",X"E6",
		X"03",X"18",X"ED",X"3A",X"84",X"4C",X"E6",X"07",X"18",X"E6",X"C9",X"C9",X"C9",X"C9",X"C9",X"C9",
		X"C9",X"C9",X"C9",X"C9",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"DD",X"77",X"06",X"23",
		X"7E",X"DD",X"77",X"07",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",X"75",X"06",
		X"DD",X"74",X"07",X"DD",X"77",X"03",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",X"23",X"DD",
		X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"04",X"C9",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"7E",
		X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"09",X"C9",X"DD",X"6E",X"06",X"DD",X"66",
		X"07",X"7E",X"23",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"77",X"0B",X"C9",X"DD",X"7E",X"02",
		X"2F",X"DD",X"A6",X"00",X"DD",X"77",X"00",X"C3",X"F4",X"2D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"4C",
		X"21",X"00",X"00",X"01",X"00",X"10",X"32",X"C0",X"50",X"79",X"86",X"4F",X"7D",X"C6",X"02",X"6F",
		X"FE",X"02",X"D2",X"09",X"30",X"24",X"10",X"EE",X"79",X"A7",X"20",X"15",X"32",X"07",X"50",X"7C",
		X"FE",X"30",X"C2",X"03",X"30",X"26",X"00",X"2C",X"7D",X"FE",X"02",X"DA",X"03",X"30",X"C3",X"42",
		X"30",X"25",X"7C",X"E6",X"F0",X"32",X"07",X"50",X"0F",X"0F",X"0F",X"0F",X"5F",X"06",X"00",X"C3",
		X"BD",X"30",X"31",X"54",X"31",X"06",X"FF",X"E1",X"D1",X"48",X"32",X"C0",X"50",X"79",X"A3",X"77",
		X"C6",X"33",X"4F",X"2C",X"7D",X"E6",X"0F",X"C2",X"4D",X"30",X"79",X"87",X"87",X"81",X"C6",X"31",
		X"4F",X"7D",X"A7",X"C2",X"4D",X"30",X"24",X"15",X"C2",X"4A",X"30",X"3B",X"3B",X"3B",X"3B",X"E1",
		X"D1",X"48",X"32",X"C0",X"50",X"79",X"A3",X"4F",X"7E",X"A3",X"B9",X"C2",X"B5",X"30",X"C6",X"33",
		X"4F",X"2C",X"7D",X"E6",X"0F",X"C2",X"75",X"30",X"79",X"87",X"87",X"81",X"C6",X"31",X"4F",X"7D",
		X"A7",X"C2",X"75",X"30",X"24",X"15",X"C2",X"72",X"30",X"3B",X"3B",X"3B",X"3B",X"78",X"D6",X"10",
		X"47",X"10",X"A4",X"F1",X"D1",X"FE",X"44",X"C2",X"45",X"30",X"7B",X"EE",X"F0",X"C2",X"45",X"30",
		X"06",X"01",X"C3",X"BD",X"30",X"7B",X"E6",X"01",X"EE",X"01",X"5F",X"06",X"00",X"31",X"C0",X"4F",
		X"D9",X"21",X"00",X"4C",X"06",X"04",X"32",X"C0",X"50",X"36",X"00",X"2C",X"20",X"FB",X"24",X"10",
		X"F5",X"21",X"00",X"40",X"06",X"04",X"32",X"C0",X"50",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",
		X"10",X"F4",X"06",X"04",X"32",X"C0",X"50",X"3E",X"0F",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F4",
		X"D9",X"10",X"08",X"06",X"23",X"CD",X"5E",X"2C",X"C3",X"74",X"31",X"7B",X"C6",X"30",X"32",X"84",
		X"41",X"C5",X"E5",X"06",X"24",X"CD",X"5E",X"2C",X"E1",X"7C",X"FE",X"40",X"2A",X"6C",X"31",X"38",
		X"11",X"FE",X"4C",X"2A",X"6E",X"31",X"30",X"0A",X"FE",X"44",X"2A",X"70",X"31",X"38",X"03",X"2A",
		X"72",X"31",X"7D",X"32",X"04",X"42",X"7C",X"32",X"64",X"42",X"3A",X"00",X"50",X"47",X"3A",X"40",
		X"50",X"B0",X"E6",X"01",X"20",X"11",X"C1",X"79",X"E6",X"0F",X"47",X"79",X"E6",X"F0",X"0F",X"0F",
		X"0F",X"0F",X"4F",X"ED",X"43",X"85",X"41",X"32",X"C0",X"50",X"3A",X"40",X"50",X"E6",X"10",X"28",
		X"F6",X"C3",X"0B",X"23",X"00",X"4C",X"0F",X"04",X"00",X"4C",X"F0",X"04",X"00",X"40",X"0F",X"04",
		X"00",X"40",X"F0",X"04",X"00",X"44",X"0F",X"04",X"00",X"44",X"F0",X"04",X"4F",X"40",X"41",X"57",
		X"41",X"56",X"41",X"43",X"21",X"06",X"50",X"3E",X"01",X"77",X"2D",X"20",X"FC",X"AF",X"32",X"03",
		X"50",X"D6",X"04",X"D3",X"00",X"31",X"C0",X"4F",X"32",X"C0",X"50",X"AF",X"32",X"00",X"4E",X"3C",
		X"32",X"01",X"4E",X"32",X"00",X"50",X"FB",X"3A",X"00",X"50",X"2F",X"47",X"E6",X"E0",X"28",X"05",
		X"3E",X"02",X"32",X"9C",X"4E",X"3A",X"40",X"50",X"2F",X"4F",X"E6",X"60",X"28",X"05",X"3E",X"01",
		X"32",X"9C",X"4E",X"78",X"B1",X"E6",X"01",X"28",X"05",X"3E",X"08",X"32",X"BC",X"4E",X"78",X"B1",
		X"E6",X"02",X"28",X"05",X"3E",X"04",X"32",X"BC",X"4E",X"78",X"B1",X"E6",X"04",X"28",X"05",X"3E",
		X"10",X"32",X"BC",X"4E",X"78",X"B1",X"E6",X"08",X"28",X"05",X"3E",X"20",X"32",X"BC",X"4E",X"3A",
		X"80",X"50",X"E6",X"03",X"C6",X"25",X"47",X"CD",X"5E",X"2C",X"3A",X"80",X"50",X"0F",X"0F",X"0F",
		X"0F",X"E6",X"03",X"FE",X"03",X"20",X"08",X"06",X"2A",X"CD",X"5E",X"2C",X"C3",X"1C",X"32",X"07",
		X"5F",X"D5",X"06",X"2B",X"CD",X"5E",X"2C",X"06",X"2E",X"CD",X"5E",X"2C",X"D1",X"16",X"00",X"21",
		X"F9",X"32",X"19",X"7E",X"32",X"2A",X"42",X"23",X"7E",X"32",X"4A",X"42",X"3A",X"80",X"50",X"0F",
		X"0F",X"E6",X"03",X"C6",X"31",X"FE",X"34",X"20",X"01",X"3C",X"32",X"0C",X"42",X"06",X"29",X"CD",
		X"5E",X"2C",X"3A",X"40",X"50",X"07",X"E6",X"01",X"C6",X"2C",X"47",X"CD",X"5E",X"2C",X"3A",X"40",
		X"50",X"E6",X"10",X"CA",X"88",X"31",X"AF",X"32",X"00",X"50",X"F3",X"21",X"07",X"50",X"AF",X"77",
		X"2D",X"20",X"FC",X"31",X"E2",X"3A",X"06",X"03",X"D9",X"E1",X"D1",X"32",X"C0",X"50",X"C1",X"3E",
		X"3C",X"77",X"23",X"72",X"23",X"10",X"F8",X"3B",X"3B",X"C1",X"71",X"23",X"3E",X"3F",X"77",X"23",
		X"10",X"F8",X"3B",X"3B",X"1D",X"C2",X"5B",X"32",X"F1",X"D9",X"10",X"DC",X"31",X"C0",X"4F",X"06",
		X"08",X"CD",X"ED",X"32",X"10",X"FB",X"32",X"C0",X"50",X"3A",X"40",X"50",X"E6",X"10",X"28",X"F6",
		X"3A",X"40",X"50",X"E6",X"60",X"C2",X"4B",X"23",X"06",X"08",X"CD",X"ED",X"32",X"10",X"FB",X"3A",
		X"40",X"50",X"E6",X"10",X"C2",X"4B",X"23",X"1E",X"01",X"06",X"04",X"32",X"C0",X"50",X"CD",X"ED",
		X"32",X"3A",X"00",X"50",X"A3",X"20",X"F4",X"CD",X"ED",X"32",X"32",X"C0",X"50",X"3A",X"00",X"50",
		X"EE",X"FF",X"20",X"F3",X"10",X"E5",X"CB",X"03",X"7B",X"FE",X"10",X"DA",X"A9",X"32",X"21",X"00",
		X"40",X"06",X"04",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F7",X"CD",X"F4",X"3A",X"32",
		X"C0",X"50",X"3A",X"40",X"50",X"E6",X"10",X"CA",X"DF",X"32",X"C3",X"4B",X"23",X"32",X"C0",X"50",
		X"21",X"00",X"28",X"2B",X"7C",X"B5",X"20",X"FB",X"C9",X"30",X"31",X"35",X"31",X"30",X"32",X"00",
		X"FF",X"01",X"00",X"00",X"01",X"FF",X"00",X"00",X"FF",X"01",X"00",X"00",X"01",X"FF",X"00",X"55",
		X"2A",X"55",X"2A",X"55",X"55",X"55",X"55",X"55",X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"25",
		X"25",X"25",X"25",X"22",X"22",X"22",X"22",X"01",X"01",X"01",X"01",X"58",X"02",X"08",X"07",X"60",
		X"09",X"10",X"0E",X"68",X"10",X"70",X"17",X"14",X"19",X"52",X"4A",X"A5",X"94",X"AA",X"2A",X"55",
		X"55",X"55",X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"92",X"24",X"25",X"49",X"48",X"24",X"22",
		X"91",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"2A",X"55",X"2A",X"55",X"55",X"55",X"55",X"AA",X"2A",X"55",X"55",X"55",
		X"2A",X"55",X"2A",X"52",X"4A",X"A5",X"94",X"48",X"24",X"22",X"91",X"21",X"44",X"44",X"08",X"58",
		X"02",X"34",X"08",X"D8",X"09",X"B4",X"0F",X"58",X"11",X"08",X"16",X"34",X"17",X"55",X"55",X"55",
		X"55",X"D5",X"6A",X"D5",X"6A",X"AA",X"6A",X"55",X"D5",X"55",X"55",X"55",X"55",X"AA",X"2A",X"55",
		X"55",X"92",X"24",X"92",X"24",X"22",X"22",X"22",X"22",X"A4",X"01",X"54",X"06",X"F8",X"07",X"A8",
		X"0C",X"D4",X"0D",X"84",X"12",X"B0",X"13",X"D5",X"6A",X"D5",X"6A",X"D6",X"5A",X"AD",X"B5",X"D6",
		X"5A",X"AD",X"B5",X"D5",X"6A",X"D5",X"6A",X"AA",X"6A",X"55",X"D5",X"92",X"24",X"25",X"49",X"48",
		X"24",X"22",X"91",X"A4",X"01",X"54",X"06",X"F8",X"07",X"A8",X"0C",X"D4",X"0D",X"FE",X"FF",X"FF",
		X"FF",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"6D",X"B6",X"6D",X"6D",X"DB",X"6D",X"6D",X"6D",
		X"6D",X"D6",X"5A",X"AD",X"B5",X"25",X"25",X"25",X"25",X"92",X"24",X"92",X"24",X"2C",X"01",X"DC",
		X"05",X"08",X"07",X"B8",X"0B",X"E4",X"0C",X"FE",X"FF",X"FF",X"FF",X"D5",X"6A",X"D5",X"6A",X"D5",
		X"6A",X"D5",X"6A",X"B6",X"6D",X"6D",X"DB",X"6D",X"6D",X"6D",X"6D",X"D6",X"5A",X"AD",X"B5",X"48",
		X"24",X"22",X"91",X"92",X"24",X"92",X"24",X"2C",X"01",X"DC",X"05",X"08",X"07",X"B8",X"0B",X"E4",
		X"0C",X"FE",X"FF",X"FF",X"FF",X"40",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",X"D2",
		X"D4",X"FC",X"FC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"D0",X"D2",X"D2",X"D2",X"D2",X"D6",
		X"D8",X"D2",X"D2",X"D2",X"D2",X"D4",X"FC",X"DA",X"09",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DC",
		X"FC",X"FC",X"FC",X"DA",X"05",X"DE",X"E4",X"05",X"DC",X"FC",X"DA",X"02",X"E6",X"E8",X"EA",X"02",
		X"E6",X"EA",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"E6",
		X"EA",X"02",X"E7",X"EB",X"02",X"E6",X"EA",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"FC",X"E4",X"02",
		X"DE",X"E4",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",
		X"E4",X"05",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"DE",X"FC",X"E4",X"02",X"DE",X"E4",X"02",
		X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"F2",X"E8",X"E8",
		X"EA",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",X"E7",X"E9",X"EB",X"02",X"E7",X"EB",X"02",
		X"E7",X"D2",X"D2",X"D2",X"EB",X"02",X"E7",X"D2",X"D2",X"D2",X"EB",X"02",X"E7",X"E9",X"E9",X"E9",
		X"EB",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"1B",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",X"02",
		X"E6",X"E8",X"F8",X"02",X"F6",X"E8",X"E8",X"E8",X"E8",X"E8",X"E8",X"F8",X"02",X"F6",X"E8",X"E8",
		X"E8",X"EA",X"02",X"E6",X"F8",X"02",X"F6",X"E8",X"E8",X"F4",X"E4",X"02",X"DC",X"FC",X"DA",X"02",
		X"DE",X"FC",X"E4",X"02",X"F7",X"E9",X"E9",X"F5",X"F3",X"E9",X"E9",X"F9",X"02",X"F7",X"E9",X"E9",
		X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"F7",X"E9",X"E9",X"F5",X"E4",X"02",X"DC",X"FC",X"DA",X"02",
		X"DE",X"FC",X"E4",X"05",X"DE",X"E4",X"0B",X"DE",X"E4",X"05",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",
		X"02",X"DE",X"FC",X"E4",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"EC",X"D3",X"D3",X"D3",X"EE",
		X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"E6",X"EA",X"02",X"DE",X"E4",X"02",X"DC",X"FC",X"DA",
		X"02",X"E7",X"E9",X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"FC",X"FC",X"DA",
		X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DE",X"E4",X"02",X"E7",X"EB",X"02",X"DC",X"FC",X"DA",
		X"06",X"DE",X"E4",X"05",X"F0",X"FC",X"FC",X"FC",X"DA",X"02",X"DE",X"E4",X"05",X"DE",X"E4",X"05",
		X"DC",X"FC",X"FA",X"E8",X"E8",X"E8",X"EA",X"02",X"DE",X"F2",X"E8",X"E8",X"EA",X"02",X"CE",X"FC",
		X"FC",X"FC",X"DA",X"02",X"DE",X"F2",X"E8",X"E8",X"EA",X"02",X"DE",X"F2",X"E8",X"E8",X"EA",X"02",
		X"DC",X"00",X"00",X"00",X"00",X"62",X"01",X"02",X"01",X"01",X"01",X"01",X"0C",X"01",X"01",X"04",
		X"01",X"01",X"01",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"04",X"03",X"0C",X"03",X"01",
		X"01",X"01",X"03",X"04",X"04",X"03",X"0C",X"06",X"03",X"04",X"04",X"03",X"0C",X"06",X"03",X"04",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",X"04",
		X"04",X"0F",X"03",X"06",X"04",X"04",X"01",X"01",X"01",X"0C",X"03",X"01",X"01",X"01",X"03",X"04",
		X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"01",X"01",
		X"01",X"01",X"03",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"08",X"18",X"08",X"18",X"04",
		X"01",X"01",X"01",X"01",X"03",X"0C",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"04",X"04",X"03",
		X"0C",X"03",X"03",X"03",X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"04",X"01",X"01",X"01",
		X"0C",X"03",X"01",X"01",X"01",X"03",X"04",X"04",X"0F",X"03",X"06",X"04",X"04",X"0F",X"03",X"06",
		X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"03",X"04",X"04",X"03",X"0C",X"06",
		X"03",X"04",X"04",X"03",X"0C",X"06",X"03",X"04",X"04",X"03",X"0C",X"03",X"01",X"01",X"01",X"03",
		X"04",X"04",X"03",X"0C",X"03",X"03",X"03",X"04",X"01",X"02",X"01",X"01",X"01",X"01",X"0C",X"01",
		X"01",X"04",X"01",X"01",X"01",X"13",X"37",X"23",X"37",X"32",X"37",X"41",X"37",X"5A",X"37",X"6A",
		X"37",X"7A",X"37",X"86",X"37",X"9D",X"37",X"B1",X"37",X"00",X"3D",X"21",X"3D",X"FD",X"37",X"67",
		X"3D",X"E3",X"3D",X"86",X"3D",X"02",X"3E",X"4C",X"38",X"5A",X"38",X"3C",X"3D",X"57",X"3D",X"D3",
		X"3D",X"76",X"3D",X"F2",X"3D",X"01",X"00",X"02",X"00",X"03",X"00",X"BC",X"38",X"C4",X"38",X"CE",
		X"38",X"D8",X"38",X"E2",X"38",X"EC",X"38",X"F6",X"38",X"00",X"39",X"0A",X"39",X"1A",X"39",X"6F",
		X"39",X"2A",X"39",X"58",X"39",X"41",X"39",X"4F",X"3E",X"86",X"39",X"97",X"39",X"B0",X"39",X"BD",
		X"39",X"CA",X"39",X"A5",X"3D",X"21",X"3E",X"C4",X"3D",X"40",X"3E",X"95",X"3D",X"11",X"3E",X"B4",
		X"3D",X"30",X"3E",X"D4",X"83",X"48",X"49",X"47",X"48",X"40",X"53",X"43",X"4F",X"52",X"45",X"2F",
		X"8F",X"2F",X"80",X"3B",X"80",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"40",X"40",X"2F",X"8F",
		X"2F",X"80",X"3B",X"80",X"46",X"52",X"45",X"45",X"40",X"50",X"4C",X"41",X"59",X"2F",X"8F",X"2F",
		X"80",X"8C",X"02",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"45",X"2F",X"85",X"2F",
		X"10",X"10",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"10",X"10",X"8C",X"02",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"40",X"54",X"57",X"4F",X"2F",X"85",X"2F",X"80",X"92",X"02",X"47",X"41",X"4D",X"45",
		X"40",X"40",X"4F",X"56",X"45",X"52",X"2F",X"81",X"2F",X"80",X"52",X"02",X"52",X"45",X"41",X"44",
		X"59",X"5B",X"2F",X"89",X"2F",X"90",X"EE",X"02",X"50",X"55",X"53",X"48",X"40",X"53",X"54",X"41",
		X"52",X"54",X"40",X"42",X"55",X"54",X"54",X"4F",X"4E",X"2F",X"87",X"2F",X"80",X"B2",X"02",X"31",
		X"40",X"50",X"4C",X"41",X"59",X"45",X"52",X"40",X"4F",X"4E",X"4C",X"59",X"40",X"2F",X"85",X"2F",
		X"80",X"B2",X"02",X"31",X"40",X"4F",X"52",X"40",X"32",X"40",X"50",X"4C",X"41",X"59",X"45",X"52",
		X"53",X"2F",X"85",X"00",X"2F",X"00",X"80",X"00",X"96",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",
		X"50",X"55",X"43",X"4B",X"4D",X"41",X"4E",X"40",X"46",X"4F",X"52",X"40",X"40",X"40",X"30",X"30",
		X"30",X"40",X"5D",X"5E",X"5F",X"2F",X"8E",X"2F",X"80",X"BA",X"02",X"5C",X"40",X"28",X"29",X"2A",
		X"2B",X"2C",X"2D",X"2E",X"40",X"31",X"39",X"38",X"30",X"2F",X"83",X"2F",X"80",X"C3",X"02",X"43",
		X"48",X"41",X"52",X"41",X"43",X"54",X"45",X"52",X"40",X"3A",X"40",X"4E",X"49",X"43",X"4B",X"4E",
		X"41",X"4D",X"45",X"2F",X"8F",X"2F",X"80",X"65",X"01",X"26",X"41",X"4B",X"41",X"42",X"45",X"49",
		X"26",X"2F",X"81",X"2F",X"80",X"45",X"01",X"26",X"4D",X"41",X"43",X"4B",X"59",X"26",X"2F",X"81",
		X"2F",X"80",X"48",X"01",X"26",X"50",X"49",X"4E",X"4B",X"59",X"26",X"2F",X"83",X"2F",X"80",X"48",
		X"01",X"26",X"4D",X"49",X"43",X"4B",X"59",X"26",X"2F",X"83",X"2F",X"80",X"76",X"02",X"10",X"40",
		X"31",X"30",X"40",X"5D",X"5E",X"5F",X"2F",X"9F",X"2F",X"80",X"78",X"02",X"14",X"40",X"35",X"30",
		X"40",X"5D",X"5E",X"5F",X"2F",X"9F",X"2F",X"80",X"5D",X"02",X"28",X"29",X"2A",X"2B",X"2C",X"2D",
		X"2E",X"2F",X"83",X"2F",X"80",X"C5",X"02",X"40",X"4F",X"49",X"4B",X"41",X"4B",X"45",X"3B",X"3B",
		X"3B",X"3B",X"2F",X"81",X"2F",X"80",X"C5",X"02",X"40",X"55",X"52",X"43",X"48",X"49",X"4E",X"3B",
		X"3B",X"3B",X"3B",X"3B",X"2F",X"81",X"2F",X"80",X"C8",X"02",X"40",X"4D",X"41",X"43",X"48",X"49",
		X"42",X"55",X"53",X"45",X"3B",X"3B",X"2F",X"83",X"2F",X"80",X"C8",X"02",X"40",X"52",X"4F",X"4D",
		X"50",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"2F",X"83",X"2F",X"80",X"12",X"02",X"81",X"85",
		X"2F",X"83",X"2F",X"90",X"32",X"02",X"40",X"82",X"85",X"40",X"2F",X"83",X"2F",X"90",X"32",X"02",
		X"40",X"83",X"85",X"40",X"2F",X"83",X"2F",X"90",X"32",X"02",X"40",X"84",X"85",X"40",X"2F",X"83",
		X"2F",X"90",X"32",X"02",X"40",X"86",X"8D",X"8E",X"2F",X"83",X"2F",X"90",X"32",X"02",X"87",X"88",
		X"8D",X"8E",X"2F",X"83",X"2F",X"90",X"32",X"02",X"89",X"8A",X"8D",X"8E",X"2F",X"83",X"2F",X"90",
		X"32",X"02",X"8B",X"8C",X"8D",X"8E",X"2F",X"83",X"2F",X"90",X"04",X"03",X"4D",X"45",X"4D",X"4F",
		X"52",X"59",X"40",X"40",X"4F",X"4B",X"2F",X"8F",X"2F",X"80",X"04",X"03",X"42",X"41",X"44",X"40",
		X"40",X"40",X"40",X"52",X"40",X"4D",X"2F",X"8F",X"2F",X"80",X"08",X"03",X"31",X"40",X"43",X"4F",
		X"49",X"4E",X"40",X"40",X"31",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"40",X"2F",X"8F",X"2F",
		X"80",X"08",X"03",X"32",X"40",X"43",X"4F",X"49",X"4E",X"53",X"40",X"31",X"40",X"43",X"52",X"45",
		X"44",X"49",X"54",X"40",X"2F",X"8F",X"2F",X"80",X"08",X"03",X"31",X"40",X"43",X"4F",X"49",X"4E",
		X"40",X"40",X"32",X"40",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"2F",X"8F",X"2F",X"80",X"08",
		X"03",X"46",X"52",X"45",X"45",X"40",X"40",X"50",X"4C",X"41",X"59",X"40",X"40",X"40",X"40",X"40",
		X"40",X"40",X"2F",X"8F",X"2F",X"80",X"0A",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"40",X"4E",
		X"4F",X"4E",X"45",X"2F",X"8F",X"2F",X"80",X"0A",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"2F",
		X"8F",X"2F",X"80",X"0C",X"03",X"50",X"55",X"43",X"4B",X"4D",X"41",X"4E",X"2F",X"8F",X"2F",X"80",
		X"0E",X"03",X"54",X"41",X"42",X"4C",X"45",X"40",X"40",X"2F",X"8F",X"2F",X"80",X"0E",X"03",X"55",
		X"50",X"52",X"49",X"47",X"48",X"54",X"2F",X"8F",X"2F",X"80",X"0A",X"02",X"30",X"30",X"30",X"2F",
		X"8F",X"2F",X"80",X"6B",X"01",X"26",X"41",X"4F",X"53",X"55",X"4B",X"45",X"26",X"2F",X"85",X"2F",
		X"80",X"4B",X"01",X"26",X"4D",X"55",X"43",X"4B",X"59",X"26",X"2F",X"85",X"2F",X"80",X"6E",X"01",
		X"26",X"47",X"55",X"5A",X"55",X"54",X"41",X"26",X"2F",X"87",X"2F",X"80",X"4E",X"01",X"26",X"4D",
		X"4F",X"43",X"4B",X"59",X"26",X"2F",X"87",X"2F",X"80",X"CB",X"02",X"40",X"4B",X"49",X"4D",X"41",
		X"47",X"55",X"52",X"45",X"3B",X"3B",X"2F",X"85",X"2F",X"80",X"CB",X"02",X"40",X"53",X"54",X"59",
		X"4C",X"49",X"53",X"54",X"3B",X"3B",X"3B",X"3B",X"2F",X"85",X"2F",X"80",X"CE",X"02",X"40",X"4F",
		X"54",X"4F",X"42",X"4F",X"4B",X"45",X"3B",X"3B",X"3B",X"2F",X"87",X"2F",X"80",X"CE",X"02",X"40",
		X"43",X"52",X"59",X"42",X"41",X"42",X"59",X"3B",X"3B",X"3B",X"3B",X"2F",X"87",X"2F",X"80",X"01",
		X"01",X"03",X"01",X"01",X"01",X"03",X"02",X"02",X"02",X"01",X"01",X"01",X"01",X"02",X"04",X"04",
		X"04",X"06",X"02",X"02",X"02",X"02",X"04",X"02",X"04",X"04",X"04",X"06",X"02",X"02",X"02",X"02",
		X"01",X"01",X"01",X"01",X"02",X"04",X"04",X"04",X"06",X"02",X"02",X"02",X"02",X"06",X"04",X"05",
		X"01",X"01",X"03",X"01",X"01",X"01",X"04",X"01",X"01",X"01",X"03",X"01",X"01",X"04",X"01",X"01",
		X"01",X"6C",X"05",X"01",X"01",X"01",X"18",X"04",X"04",X"18",X"05",X"01",X"01",X"01",X"17",X"02",
		X"03",X"04",X"16",X"04",X"03",X"01",X"01",X"01",X"76",X"01",X"01",X"01",X"01",X"03",X"01",X"01",
		X"01",X"02",X"04",X"02",X"04",X"0E",X"02",X"04",X"02",X"04",X"02",X"04",X"0B",X"01",X"01",X"01",
		X"02",X"04",X"02",X"01",X"01",X"01",X"01",X"02",X"02",X"02",X"0E",X"02",X"04",X"02",X"04",X"02",
		X"01",X"02",X"01",X"0A",X"01",X"01",X"01",X"01",X"03",X"01",X"01",X"01",X"03",X"01",X"01",X"03",
		X"04",X"00",X"02",X"40",X"01",X"3E",X"3D",X"10",X"40",X"40",X"0E",X"3D",X"3E",X"10",X"C2",X"43",
		X"01",X"3E",X"3D",X"10",X"21",X"A2",X"40",X"11",X"4F",X"3A",X"36",X"14",X"1A",X"A7",X"C8",X"13",
		X"85",X"6F",X"D2",X"FA",X"3A",X"24",X"18",X"F2",X"90",X"14",X"94",X"0F",X"98",X"15",X"98",X"15",
		X"A0",X"14",X"A0",X"14",X"A4",X"17",X"A4",X"17",X"A8",X"09",X"A8",X"09",X"9C",X"16",X"9C",X"16",
		X"AC",X"16",X"AC",X"16",X"AC",X"16",X"AC",X"16",X"AC",X"16",X"AC",X"16",X"AC",X"16",X"AC",X"16",
		X"73",X"20",X"00",X"0C",X"00",X"0A",X"1F",X"00",X"72",X"20",X"FB",X"87",X"00",X"02",X"0F",X"00",
		X"36",X"20",X"04",X"8C",X"00",X"00",X"06",X"00",X"36",X"28",X"05",X"8B",X"00",X"00",X"06",X"00",
		X"36",X"30",X"06",X"8A",X"00",X"00",X"06",X"00",X"36",X"3C",X"07",X"89",X"00",X"00",X"06",X"00",
		X"36",X"48",X"08",X"88",X"00",X"00",X"06",X"00",X"24",X"00",X"06",X"08",X"00",X"00",X"0A",X"00",
		X"40",X"70",X"FA",X"10",X"00",X"00",X"0A",X"00",X"70",X"04",X"00",X"00",X"00",X"00",X"08",X"00",
		X"42",X"18",X"FD",X"06",X"00",X"01",X"0C",X"00",X"42",X"04",X"03",X"06",X"00",X"01",X"0C",X"00",
		X"56",X"0C",X"FF",X"8C",X"00",X"02",X"0F",X"00",X"05",X"00",X"02",X"20",X"00",X"01",X"0C",X"00",
		X"41",X"20",X"FF",X"86",X"FE",X"1C",X"0F",X"FF",X"70",X"00",X"01",X"0C",X"00",X"01",X"08",X"00",
		X"01",X"02",X"04",X"08",X"10",X"20",X"40",X"80",X"00",X"57",X"5C",X"61",X"67",X"6D",X"74",X"7B",
		X"82",X"8A",X"92",X"9A",X"A3",X"AD",X"B8",X"C3",X"D4",X"3B",X"F3",X"3B",X"58",X"3C",X"95",X"3C",
		X"DE",X"3C",X"DF",X"3C",X"F1",X"02",X"F2",X"03",X"F3",X"0F",X"F4",X"01",X"82",X"70",X"69",X"82",
		X"70",X"69",X"83",X"70",X"6A",X"83",X"70",X"6A",X"82",X"70",X"69",X"82",X"70",X"69",X"89",X"8B",
		X"8D",X"8E",X"FF",X"F1",X"02",X"F2",X"03",X"F3",X"0F",X"F4",X"01",X"67",X"50",X"30",X"47",X"30",
		X"67",X"50",X"30",X"47",X"30",X"67",X"50",X"30",X"47",X"30",X"4B",X"10",X"4C",X"10",X"4D",X"10",
		X"4E",X"10",X"67",X"50",X"30",X"47",X"30",X"67",X"50",X"30",X"47",X"30",X"67",X"50",X"30",X"47",
		X"30",X"4B",X"10",X"4C",X"10",X"4D",X"10",X"4E",X"10",X"67",X"50",X"30",X"47",X"30",X"67",X"50",
		X"30",X"47",X"30",X"67",X"50",X"30",X"47",X"30",X"4B",X"10",X"4C",X"10",X"4D",X"10",X"4E",X"10",
		X"77",X"20",X"4E",X"10",X"4D",X"10",X"4C",X"10",X"4A",X"10",X"47",X"10",X"46",X"10",X"65",X"30",
		X"66",X"30",X"67",X"40",X"70",X"F0",X"FB",X"3B",X"F1",X"00",X"F2",X"02",X"F3",X"0F",X"F4",X"00",
		X"42",X"50",X"4E",X"50",X"49",X"50",X"46",X"50",X"4E",X"49",X"70",X"66",X"70",X"43",X"50",X"4F",
		X"50",X"4A",X"50",X"47",X"50",X"4F",X"4A",X"70",X"67",X"70",X"42",X"50",X"4E",X"50",X"49",X"50",
		X"46",X"50",X"4E",X"49",X"70",X"66",X"70",X"45",X"46",X"47",X"50",X"47",X"48",X"49",X"50",X"49",
		X"4A",X"4B",X"50",X"6E",X"FF",X"F1",X"01",X"F2",X"01",X"F3",X"0F",X"F4",X"00",X"26",X"67",X"26",
		X"67",X"26",X"67",X"23",X"44",X"42",X"47",X"30",X"67",X"2A",X"8B",X"70",X"26",X"67",X"26",X"67",
		X"26",X"67",X"23",X"44",X"42",X"47",X"30",X"67",X"23",X"84",X"70",X"26",X"67",X"26",X"67",X"26",
		X"67",X"23",X"44",X"42",X"47",X"30",X"67",X"29",X"6A",X"2B",X"6C",X"30",X"2C",X"6D",X"40",X"2B",
		X"6C",X"29",X"6A",X"67",X"20",X"29",X"6A",X"40",X"26",X"87",X"70",X"F0",X"9D",X"3C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"03",X"42",X"4F",X"4E",X"55",X"53",X"40",X"50",X"41",X"43",X"3B",X"4D",X"41",X"4E",X"40",
		X"46",X"4F",X"52",X"40",X"40",X"40",X"30",X"30",X"30",X"40",X"5D",X"5E",X"5F",X"2F",X"8E",X"2F",
		X"80",X"3A",X"03",X"5C",X"40",X"31",X"39",X"38",X"30",X"40",X"4D",X"49",X"44",X"57",X"41",X"59",
		X"40",X"4D",X"46",X"47",X"25",X"43",X"4F",X"25",X"2F",X"83",X"2F",X"80",X"3D",X"03",X"5C",X"40",
		X"31",X"39",X"38",X"30",X"40",X"4D",X"49",X"44",X"57",X"41",X"59",X"40",X"4D",X"46",X"47",X"25",
		X"43",X"4F",X"25",X"2F",X"83",X"2F",X"80",X"C5",X"02",X"3B",X"53",X"48",X"41",X"44",X"4F",X"57",
		X"40",X"40",X"40",X"2F",X"81",X"2F",X"80",X"65",X"01",X"26",X"42",X"4C",X"49",X"4E",X"4B",X"59",
		X"26",X"40",X"2F",X"81",X"2F",X"80",X"C8",X"02",X"3B",X"53",X"50",X"45",X"45",X"44",X"59",X"40",
		X"40",X"40",X"2F",X"83",X"2F",X"80",X"68",X"01",X"26",X"50",X"49",X"4E",X"4B",X"59",X"26",X"40",
		X"40",X"2F",X"83",X"2F",X"80",X"CB",X"02",X"3B",X"42",X"41",X"53",X"48",X"46",X"55",X"4C",X"40",
		X"40",X"2F",X"85",X"2F",X"80",X"6B",X"01",X"26",X"49",X"4E",X"4B",X"59",X"26",X"40",X"40",X"40",
		X"2F",X"85",X"2F",X"80",X"CE",X"02",X"3B",X"50",X"4F",X"4B",X"45",X"59",X"40",X"40",X"40",X"40",
		X"2F",X"87",X"2F",X"80",X"6E",X"01",X"26",X"43",X"4C",X"59",X"44",X"45",X"26",X"40",X"40",X"2F",
		X"87",X"2F",X"80",X"C5",X"02",X"3B",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"41",X"3B",X"2F",
		X"81",X"2F",X"80",X"65",X"01",X"26",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"26",X"2F",X"81",
		X"2F",X"80",X"C8",X"02",X"3B",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"43",X"3B",X"2F",X"83",
		X"2F",X"80",X"68",X"01",X"26",X"44",X"44",X"44",X"44",X"44",X"44",X"44",X"26",X"2F",X"83",X"2F",
		X"80",X"CB",X"02",X"3B",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"45",X"3B",X"2F",X"85",X"2F",
		X"80",X"6B",X"01",X"26",X"46",X"46",X"46",X"46",X"46",X"46",X"46",X"26",X"2F",X"85",X"2F",X"80",
		X"CE",X"02",X"3B",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"47",X"3B",X"2F",X"87",X"2F",X"80",
		X"6E",X"01",X"26",X"48",X"48",X"48",X"48",X"48",X"48",X"48",X"26",X"2F",X"87",X"2F",X"80",X"0C",
		X"03",X"50",X"41",X"43",X"3B",X"4D",X"41",X"4E",X"2F",X"8F",X"2F",X"80",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"8D",X"00",X"75",X"73");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
